module lut_weights_1(sbyte,addr);
input [3:0] addr;
output reg [1727:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0001: sbyte = 1728'b000000000011100000000000001010010000000000010110000000000110000000000000001001111111111111111101000000000101100100000000000010101111111111110111111111111101100100000000000100001111111111101110111111111010100111111111110000101111111110101011111111111100000111111111110101101111111110111000111111111010101111111111100100011111111111010011111111111110000111111111111000100000000000001011000000000110011100000000011000010000000001000100111111111101100011111111110011111111111111110110111111111111111100000000010001100000000001011111000000000001010000000000001110010000000001011010111111111100011111111111111000101111111111110000000000000001011100000000000001011111111111111001000000000001110100000000000111010000000000101111000000000011101000000000001101110000000000110001000000000100001000000000001101000000000000100111000000000011000100000000001100011111111111111100000000000010110100000000000100100000000000101101111111111111000111111111110110011111111111100101111111111110001111111111110101111111111111101011111111111111111000000000000000001111111111110100000000000000011000000000000000010000000000001101111111111101110011111111111111110000000000001101111111111111110011111111110001001111111111010011111111111100000100000000001001100000000000011100111111111111100000000000001100000000000000100001111111111111000011111111111101011111111111110111000000000001000011111111111101010000000000000000111111111111111000000000001011100000000000000001111111111111010100000000001100000000000000011111000000000010100000000000101001100000000001110011000000000100001100000000011011010000000001010000111111111111011011111111111100101111111110110101000000000000000100000000001101001111111111011101000000000010000100000000001011110000000000010111;
endcase
end
endmodule



module lut_weights_2(sbyte,addr);
input [3:0] addr;
output reg [20735:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0010: sbyte = 20736'b000000000000100100000000000101011111111111011101000000000001001000000000000000100000000000001111000000000000100000000000000010110000000000001110000000000000011011111111111111000000000000010101111111111111011100000000000000000000000000010001111111111111101111111111111111111111111111110110111111111111101011111111111100111111111111111111111111111101111111111111111111000000000000011011111111111110010111111111110100010000000000000001000000000000110000000000000110011111111111110110111111111111011100000000000011111111111111101111111111111111010011111111111111010000000000000010111111111111111111111111111111110000000000010101111111111111001011111111111110001111111111110001000000000001000100000000000101011111111111110100111111111111110011111111110110011111111111111000111111111111100000000000000001010000000000000000000000000000001100000000000100101111111111111101111111111111101100000000000010001111111111110010111111111110001111111111111110001111111111101110111111111111111111111111111010100000000000010010000000000000011100000000000011101111111111111111000000000001011011111111111100010000000000000010000000000010000111111111111010100000000000000111000000000000011100000000000101110000000000010010111111111111111011111111111100101111111111101111000000000010000000000000000101011111111111101110000000000001100011111111111010001111111111101101111111111111001000000000000110001111111111111011000000000000111000000000000000011111111111110101000000000000100011111111111110011111111111111111111111111101101011111111111111101111111111100101111111111110100000000000000000111111111111110111111111111111010100000000000010010000000000000100000000000000110011111111111010110000000000001011000000000000010111111111111011111111111111111010111111111111010100000000000001100000000000111110111111111101001100000000000000010000000000101000111111111101111111111111111111100000000000011000000000000000010111111111111000101111111111001111111111111111011111111111110111011111111111100101000000000010111000000000000001100000000000000000111111111111010000000000000001011111111111101110111111111110010111111111110100101111111110101100111111111110011111111111101010101111111110110100000000000001011100000000001110010000000000001011000000000011000100000000000000011111111111110110111111111101001011111111111010101111111111011101111111111100011011111111111101101111111111110001000000000000000111111111111100011111111111111000111111111101100011111111111100001111111111101101000000000000001100000000001100010000000000111000111111111111001000000000001100000000000000110010111111111101101000000000001000111111111111111011000000000000100011111111111111111111111111111010111111111111111011111111111011001111111111110000000000000001011000000000001010000000000000001010000000000001000100000000000100001111111111111110000000000000000000000000000111011111111111110010000000000000010011111111111110110000000000011111000000000000111000000000000110100000000000010101000000000010000000000000000011011111111111010000111111111110111011111111111001100000000000000101111111111111111100000000000001010000000000101001111111111111111100000000000100100000000000000010111111111110110000000000000000110000000000000101000000000001100000000000011110010000000001101010000000000000101100000000010011100000000000101011111111111100011111111111111100111111111111010110000000000000001100000000000011000000000000100100000000000000000000000000000001011111111111111101111111111101100011111111111110100000000000010010111111111110100111111111111010011111111111111100111111111110101011111111111111000000000000110001111111111111111000000000000000000000000000001111000000000001111000000000000000111111111111100010111111111111110011111111111101101111111111011011000000000001001011111111111111001111111111110001111111111110111100000000000110100000000000010111000000000001101011111111111011001111111111011111000000000000100111111111110100011111111110100110000000000000100100000000010011110000000000110110000000000000101100000000001100010000000000100001000000000001010000000000000001111111111111111100000000000000101000000000000000100000000000000001111111111111011011111111111010110000000000001001000000000001101111111111111110101111111111100111111111111111100100000000000011001111111111111110111111111110100011111111111001010000000000100010111111111110110000000000000010011111111111110000000000000001100111111111111011111111111111101000000000000000110011111111111000101111111111110001000000000001110011111111111000110000000000000110000000000000000100000000000010101111111111111111000000000001101111111111111011011111111111110010111111111111001111111111111011100000000000011110000000000001110100000000000010110000000000111100000000000011010100000000000010100000000000001111000000000000100111111111111111001111111111011110000000000000111000000000000010000000000000010110000000000001000000000000000000100000000000001111111111111111011011111111111010011111111111110110111111111110110000000000001010100000000000100100000000000000001100000000001101000000000000001011000000000001001000000000000011111111111111111001111111111111110100000000001010110000000000110110000000000000100111111111111110000000000000000110111111111111001011111111111110000000000000010111111111111110111111111111111110110000000000001011000000000000110111111111111011011111111111111011111111111111001111111111111110111111111111101001000000000001110111111111111010111111111111110110000000000000111011111111111010110000000000000000000000000001011000000000000101101111111111110111000000000001000000000000000010000000000000000101000000000000000111111111111011110000000000000011000000000000010000000000000010111111111111111011111111111111010100000000001010100000000000010001000000000000000000000000000101101111111111101000111111111111011100000000000011101111111111100111111111111111100111111111111110010000000000011100000000000000010100000000000011100000000000010010111111111111001100000000000000110000000000000110000000000000010100000000000100010000000000001001111111111111011111111111111010011111111111111000111111111110111011111111111010111111111111111111000000000010100000000000000011110000000000001000000000000001001100000000000011111111111111110111000000000000000100000000001001011111111111111110000000000000001111111111111110000000000000101001111111111111100100000000000001001111111111110110000000000001100000000000000101000000000000000000111111111111100111111111111110101111111111110100000000000000010100000000000011111111111111110111111111111111010100000000000101110000000000010110111111111110000011111111110110010000000000010110111111111111111111111111111110111111111111111000000000000001101011111111111100110000000000001010111111111110101011111111111010110000000000100110111111111111100111111111111011000000000000100001111111111111010100000000000000011111111111101111111111111111111111111111111100111111111111111000111111111111101011111111111101100000000000010001111111111111111000000000000001111111111111111010111111111111011011111111111011110000000000000111000000000001000111111111110100111111111111111100111111111111100111111111111011010000000000001011111111111111101011111111110101100000000000000000111111111110101111111111111111111111111111111010000000000001101100000000001011011111111111101111111111111111101100000000000100001111111111101110111111111110101000000000000000111111111111100110111111111111111111111111111111101111111111111010000000000000000011111111111110111111111111111000000000000000000011111111111110101111111111111010000000000000010000000000000010101111111111110101111111111111000011111111111100100000000000001111000000000000101100000000000111111111111111111111000000000001100000000000000101000000000000000110111111111111100111111111111110101111111111110010000000000000001000000000000010000000000000001001000000000000101100000000000011001111111111110100000000000001010111111111111110101111111111110101000000000001000000000000000011110000000000001011111111111111101000000000000011110000000000010001111111111111011100000000001001100000000000001001111111111111100011111111111110000000000000011000000000000000111000000000000000010000000000000100000000000001010111111111111010010000000000001001000000000001011000000000000010111111111111101110000000000000110000000000000010101111111111110001111111111110110111111111111110100000000000010100111111111111011000000000001001111111111111101111000000000000100000000000000000101111111111110110111111111111101111111111111110010000000000000000111111111110111000000000000000001111111111101101000000000001001011111111111100010000000000011100000000000000001000000000000000001111111111100001000000000000000011111111111110000000000000010001111111111110101011111111111100000000000000000110000000000000001111111111111110000000000000000101111111111110011111111111111001010000000000001111111111111111001000000000000000011111111111101010000000000000110100000000000111000000000000100000000000000001001100000000000100010000000000010010000000000010110000000000001100100000000000010111000000000001011011111111111111110000000000000001000000000000110111111111111100101111111111110110000000000000110111111111111111110000000000001001111111111110111100000000000010010000000000010010111111111110101000000000000001000000000000000100111111111110100000000000000011001111111111110110000000000001100111111111111111100000000000000010000000000001001100000000000001010000000000000010000000000000101000000000000011101111111111111010000000000000011000000000000000001111111111110001111111111110010000000000000000001111111111010101111111111111001111111111111100101111111111110100111111111111111000000000000111110000000000001011000000000010011011111111111101011111111111111011111111111111000111111111111101110000000000000110111111111111000100000000001101101111111111111110000000000000001011111111111111000000000000000001000000000001101111111111111100100000000000000100111111111111001011111111111110111111111111100110000000000001001000000000000010000000000000001010000000000010110000000000001000010000000000100010111111111110101111111111111110001111111111111101000000000000001100000000000101111111111111111101000000000010010000000000000100010000000000010110111111111111110111111111111011001111111111101110111111111110110100000000000100001111111111111111000000000000101011111111110111110000000000000110111111111111101011111111111100000000000000000101000000000000111000000000000001111111111111101100000000000000111100000000000001010000000000010110000000000001000011111111111001000000000000000011000000000001001100000000000000000000000000000011111111111111110111111111111010100000000000010110000000000000000011111111111011001111111111111110111111111110100011111111111101111111111111101111000000000001001011111111111011111111111111111011000000000001001100000000000010110000000000000000000000000000010100000000001000111111111111101001000000000001011111111111111110111111111111101101111111111110101000000000000010111111111111101010111111111110101100000000001000111111111111100011111111111111001111111111111110101111111111010010000000000000101100000000000111101111111111111110000000000000100111111111111010101111111111101010111111111111100011111111111110001111111111101010111111111101111111111111111011000000000000010001111111111111100011111111111111010000000000100100111111111111110100000000000001000000000000010100000000000000011111111111111100011111111111110001111111111111000011111111111110101111111111110000000000000001000100000000000000100000000000010001000000000000010000000000000000001111111111011011000000000001111011111111111100011111111111100110000000000001000111111111111100011111111111101001000000000000101000000000000100110000000000001101000000000000110100000000000010011111111111110011000000000000000111111111111011110000000000010011000000000000001100000000000001110000000000001000000000000000011000000000000100111111111111110101111111111111001000000000000110000000000000001111000000000000110000000000000110010000000000110100000000000000111100000000000110000000000000000110111111111111100100000000000010101111111111111100111111111111010011111111111111110000000000000111111111111111101111111111111101100000000000010000111111111111010111111111111100101111111111110101111111111111000000000000000010001111111111110111111111111110110111111111111110010000000000001111111111111110100011111111110110111111111111010100000000000000011000000000000101010000000000101100000000000000101000000000000000010000000000000111000000000010101100000000001000000000000000101110000000000000110111111111111101111111111111011110000000000000011011111111111100110000000000010010000000000001011100000000000000111111111111111101000000000001001111111111111100111111111111100110000000000001000100000000000011101111111111101011111111111110110111111111111111001111111111110001000000000000011111111111111010100000000000000010000000000000011100000000000001011111111111110001000000000000110111111111111111101111111111111110000000000000011111111111111110101111111111100110000000000000001011111111110100001111111111101001111111111110100011111111111101100000000000000111000000000000001000000000000001100000000000000000000000000001111000000000000110100000000000000001000000000000000100000000000010110000000000001000111111111111110000000000000100100000000000000111111111111111101111111111111110001111111111111110000000000000001000000000000101111111111111110111111111111111101000000000000011001111111111110000000000000000010100000000000111100000000000101010111111111110101111111111111101110000000000100110000000000001101000000000000000010000000000010101000000000000000111111111111110111111111111101010000000000000110100000000000001010000000000010111000000000000100111111111111001111111111111101001000000000001001011111111111111101111111111111011000000000000010111111111111101100000000000000010111111111111100011111111111100010000000000001011111111111111100000000000000100100000000000010000000000000000110100000000000010000000000000001011111111111111011011111111110101111111111111010111111111111110000111111111111010101111111111110100111111111110110111111111111001001111111111011010000000000011011100000000001000010000000000011011000000000010011100000000001100110000000001000000000000000010101100000000000010100000000000001101111111111111011011111111111101111111111111111011111111111110111111111111111100000000000000010010000000000011000011111111111111101111111111101110111111111110110000000000001001011111111111010011111111111110111011111111111100001111111111001100111111111110111000000000001000101111111111101000000000000010010011111111111111010000000000000100000000000000001111111111111101100000000000001111000000000000111100000000000000000000000000001010111111111101111111111111111010011111111111011011111111111101110000000000000000001111111111011001111111111111011000000000000000101111111111100100000000000000011100000000000110000000000000010111000000000000110000000000000101010000000000110000000000000001001011111111111011100000000000011011000000000000000000000000000001100000000000000101111111111111000000000000000001110000000000000100111111111110100011111111111100110000000000000000000000000010101100000000000101000000000000100111000000000000111100000000000101000000000000001111000000000001101000000000001001110000000000000111111111111111010100000000000011000000000000001110000000000000010100000000001000100000000000010111000000000000011000000000000000011111111111101111111111111111011011111111111101001111111111010101111111111110001111111111111100001111111111000100111111111110010000000000000000011111111111011001000000000001101111111111111011000000000000000111000000000000110000000000000101010000000000100111111111111111100000000000000110010000000000101111111111111110001011111111111001011111111111110000111111111110001000000000000101110000000000101111111111111111011111111111111101010000000000000011111111111111111111111111110101111111111111100111000000000001100111111111111010001111111111010110111111111110011011111111111011100000000000000011111111111101100100000000000010100000000000010111111111111111011100000000000010001111111111101110111111111111100111111111110010011111111110111010111111111111101000000000001011000000000000100001000000000011111000000000000101010000000000010111000000000001011111111111111110110000000000010100111111111110010011111111111100100000000000010001000000000000000011111111111101011111111111101111111111111111001111111111110111001111111111111000111111111101110000000000000001111111111111011110111111111110101000000000001000010000000000001111111111111111111000000000000000110000000000001100111111111111101111111111110101101111111111110101000000000000100111111111110100101111111111101000000000000001111011111111111010001111111111011011111111111110100011111111111101101111111111110110000000000000000011111111111011100000000000000111000000000001000100000000000010010000000000000011000000000010000000000000001000010000000000100110000000000100000111111111111111000000000000000110000000000001100011111111111011110000000000000011000000000000101000000000000110010000000000001100000000000000000011111111111100110000000000000000000000000001110011111111111111011111111111110001111111111111100000000000000110000000000000011000111111111111100000000000010011100000000001000010111111111111110000000000001100000000000000001101111111111111011100000000001011110000000001000010111111111111110000000000000011000000000000010100111111111111010011111111110111010000000000010010111111111111011000000000000010110000000000000001000000000000000000000000000011001111111111110111000000000000010011111111111100000000000000000000000000000000010100000000000010010000000000001100111111111111101011111111110111000000000000010001000000000000001100000000000000110000000000001100000000000000000000000000000001110000000000001010000000000001011111111111111111000000000000000000111111111101111100000000000011111111111111100010111111111110111000000000000001111111111111101111000000000001011111111111111101110000000000001111111111111110011000000000000001010000000000000001000000000000110011111111111000101111111111111101000000000000111000000000001001110000000000011100000000000000101111111111111101100000000000001110111111111110110011111111111010101111111111110000000000000000000011111111111110111111111111111010111111111111110011111111111110011111111111110110000000000000001111111111111100001111111111110010111111111110110000000000000001111111111111110110000000000000001111111111111010100000000000000001111111111110111000000000000000110000000000001001000000000000100000000000000011001111111111110000000000000000100011111111111111101111111111111110111111111111101100000000000000000000000000010000111111111111011011111111111110010000000000010010000000000000011000000000000000100000000000001111111111111111101000000000000011110000000000010111111111111111000011111111111010100000000000000000000000000001101100000000000100011111111111110111111111111111011111111111111100111111111111100011111111111111010100000000000001000000000000000101000000000001001111111111111100000000000000000110111111111111101111111111111000011111111111011110000000000001011100000000000010111111111111111000000000000010000111111111111011111111111111110011000000000000111111111111111010100000000000010010111111111110101100000000000100110000000000001111000000000001100100000000000101110000000000000010000000000000001000000000000000101111111111101001111111111111101111111111111100100000000000000110111111111111101100000000000101111111111111110011111111111110110111111111111111011111111111110010111111111111111100000000000011110000000000000100111111111111000100000000000000101111111111110010000000000001111000000000000010000000000000000001000000000001010111111111111010000000000000011011000000000001101000000000000001010000000000001110000000000000001100000000000010100000000000000011111111111111111100000000000010000000000000000010111111111110111011111111111110111111111111110001111111111111101100000000000000000000000000011010111111111111001100000000000110000000000000011001111111111110111000000000000011010000000000010010111111111101100011111111111010010000000000000011111111111111110011111111111101111111111111111010111111111111010000000000000001001111111111111000111111111111000000000000001000000000000000010001000000000000001100000000000010010000000000001011000000000000111100000000000001001111111111100111111111111101100111111111111010011111111111110011111111111110101100000000000011000000000000000101111111111111000111111111111111001111111111111010111111111101100011111111111100100000000000000000000000000000111111111111111100111111111111010101111111111111011011111111111110100000000000000010111111111110111011111111111011110000000000001101000000000000001011111111111001111111111111111101111111111110110111111111111110100000000000000100111111111111011100000000000101101111111111110111000000000000000011111111111010110000000000001111111111111111100000000000000011001111111111111001;
endcase
end
endmodule



module lut_weights_3(sbyte,addr);
input [3:0] addr;
output reg [20735:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0011: sbyte = 20736'b111111111111111100000000000100111111111111101100111111111111110100000000000000100000000000010101000000000000101100000000000001001111111111010110111111111100110111111111101101001111111110111111111111111111001000000000000100000000000000011111000000000011000000000000001000100000000000110110111111111101110000000000000001010000000000001011000000000000100000000000001000110000000000010010000000000011010000000000001001100000000000010000000000000000010100000000000011101111111111110011111111111101111011111111111011010000000000001011000000000000000000000000000100001111111111111110111111111111010000000000000011101111111111111100111111111111101111111111111100011111111111100011000000000000110000000000000101001111111111111001111111111111100100000000000010110000000000101101111111111110110111111111111110001111111111110001111111111110100111111111111011101111111111011110111111111110100111111111111101100000000000011001111111111111100000000000000010100000000000100101000000000000010000000000000101110000000000001011000000000001100100000000000010101111111111111000000000000000110111111111111101100000000000001101111111111110001111111111111011111111111111110101000000000100011100000000001010000000000000011101000000000000010100000000000001000000000000000000111111111110100000000000000000111111111111101111111111111100111011111111111011101111111111111100000000000001010000000000001101100000000000101000000000000001001000000000001000110000000000011011111111111110011111111111111110111111111111111010000000000000010000000000000000011111111111101111111111111111100100000000000010011111111111100101000000000000100100000000000001101111111111111001111111111111101100000000000010000000000000101111111111111110001011111111111101110000000000100001000000000000100100000000000000110000000000000000000000000000111000000000001010001111111111111010000000000010010000000000000111111111111111111010000000000011000100000000001001100000000000000110000000000010101000000000000011111111111111011110000000000010000011111111111110101111111111010110000000000011011000000000000110011111111111100111000000000011011111111111111001111111111111010011000000000001101011111111111010101111111111011000000000000010100000000000000100101111111111110101111111111110100111111111111101100000000000011000000000000000000011111111111001100000000000000011000000000010000100000000000110001111111111101010111111111110001000000000000000111111111111111101111111111110100011111111111111001111111111110000000000000001101011111111111000100000000000010001111111111111001011111111111100111111111111111000000000000000110100000000000010000000000000000001000000000000010100000000000110101111111111110000000000000000000000000000000010111111111111101001000000000001000011111111111111111111111111110001111111111111110000000000000011100000000000010101000000000000001100000000001000001111111111110111000000000001101100000000000011010000000000001111111111111111000000000000000101001111111111101001111111111110000100000000000001110000000000000111000000000000000011111111111010100000000000000001000000000010100000000000000010101111111111011011000000000010110111111111111010011111111111110011000000000000110011111111111110011111111111100111000000000000000011111111111010100000000000000111111111111111011111111111111011010000000000010111000000000000100011111111111111001111111111111101000000000000000000000000000001100000000000010001000000000000010100000000000000000000000000010010111111111111110000000000000110101111111111110001111111111111010000000000000010100000000000011110000000000001011011111111111111110000000000000101000000000000011000000000000001100000000000000110111111111110100100000000000100001111111111111000000000000000101011111111111011100000000000010000000000000000000000000000000100010000000000000000000000000011000011111111111100101111111111111000000000000000101111111111111011001111111111101011111111111110011100000000000011110000000000011001111111111111010100000000000000110000000000000101000000000000000111111111111110001111111111100111000000000000100111111111111000100000000000000001111111111110011011111111111110001111111111110111000000000000011100000000000011100000000000001011111111111111111000000000000000001111111111110100111111111110011011111111111100110000000000011011000000000010000111111111111101101111111111011110000000000001000111111111111110110000000000001011111111111111111011111111111111011111111111111100111111111101101111111111111101011111111111111011111111111110101100000000000011100000000000000111000000000000100100000000000101010000000000000011111111111110001111111111111101110000000000000010000000000000000111111111111100011111111111101111111111111111110000000000000001011111111111111110000000000000101100000000000000010000000000000000111111111111101111111111111101110000000000010000000000000000010011111111111101000000000000000101111111111110111011111111111111110000000000001100111111111111110100000000000010101111111111110101000000000000100000000000001010000000000000010110000000000000110111111111111011001111111111111111111111111111011111111111111110110000000000010000000000000000011000000000000010100000000000010100000000000000110000000000000000111111111111111101000000000000001000000000000110101111111111111100111111111111001011111111111111010000000000000000111111111111100011111111111110110000000000001000000000000001100111111111111100010000000000001101000000000000001000000000000010010000000000011100000000000001001100000000000110001111111111111100000000000001010100000000000101101111111111101110000000000000111000000000001001100000000000011001000000000101100100000000000100101111111111110000000000000000111111111111111011111111111111101100111111111111000000000000000011001111111111100101000000000001000100000000000011100000000000000101111111111111111100000000000111000000000000011011000000000000000100000000000100110000000000011011111111111110100100000000000010111111111111100100000000000001010011111111111100110000000000000010111111111111111011111111111111001111111111100001000000000000000100000000000010101111111111010000111111111110111111111111111111010000000000000011000000000001001100000000000000001111111111110000000000000000001000000000000001101111111111101000000000000000100011111111111001111111111111101000000000000000101000000000000000011111111111111011111111111110011111111111111111001111111111110110000000000011011011111111111111111111111111110100000000000010010011111111111101101111111111101101111111111110011000000000000001111111111111101110111111111111101111111111111101000000000000001010000000000001001100000000000110100000000000001010000000000010110000000000001010011111111111110111000000000010000011111111111101110000000000000101111111111110110100000000000000000000000000000100000000000000000011111111111110001111111111110111111111111111001000000000000000010000000000001100111111111111100100000000000100101111111111110100000000000000001111111111111011100000000000010010111111111110100111111111111110010000000000001100111111111111001100000000000011100000000000001001111111111111000111111111111101100000000000000000111111111111001100000000000001010000000000001001000000000000100000000000000110011111111111101001111111111111111111111111111110111111111111110001000000000000111011111111111110110000000000010011000000000000000000000000000000101111111111110111000000000000000011111111111011100000000000011111111111111110010011111111111100010000000000000010111111111111001111111111111110101111111111100111111111111110101000000000001000100000000000000110000000000001001011111111111101100000000000011010111111111111001111111111111101010000000000000011000000000000010000000000000000101111111111111001000000000001010100000000000101000000000000010100000000000000010100000000000000001111111111011111000000000001010111111111111011101111111111110100111111111110100111111111111101010000000000010111000000000010011111111111111010101111111111110101000000000000101100000000000100100000000000001011111111111111000111111111110111111111111111111010000000000001011000000000000001101111111111110101111111111111010111111111111011110000000000001011000000000000100111111111111101000000000000001001000000000000000011111111111100011111111111100010000000000000110000000000000010100000000000000110111111111111000111111111111100110000000000000001000000000000000111111111111101101111111111110001111111111110101011111111111000110000000000000011000000000000111100000000000110010000000000010000000000000000100111111111110111101111111111101010000000000000000000000000000101010000000000010011111111111111111100000000000001001111111111111010000000000000011000000000000001010000000000001111000000000000011100000000000000110000000000001111111111111111101100000000000001100000000000000101111111111111111011111111111101101111111111111001000000000001010111111111111110011111111111111011111111111110110011111111111111111111111111110110111111111110101100000000000001111111111111101011000000000000011100000000000101100000000000000001111111111111010100000000000000010000000000101000000000000000100000000000000000010000000000001011111111111111111100000000000111110000000000001111111111111111100100000000000100110000000000000110000000000000001100000000000001011111111111111100000000000000001011111111111010100000000000000001000000000000010000000000000010000000000000000001111111111110101000000000000011100000000000001011111111111111111111111111111001111111111111100110000000000000000100000000000100010000000000000000111111111110101111111111111110101111111111011100000000000000100100000000000100011111111111111111000000000000000000000000000000110000000000000011000000000000011111111111111100010000000000000100111111111111000011111111111110100000000000000010000000000000010000000000001010111111111111111000000000000000111100000000000100111111111111111010111111111111010011111111111011111111111111110101111111111111000100000000000010101111111111111010111111111111101011111111111111001111111111110101000000000000111011111111111111110000000000000000000000000000011011111111110111101111111111100101111111111111100000000000000101100000000000101010111111111110111000000000000111010000000000101111111111111111111100000000000011110000000000001010000000000000110111111111111010000000000000000111111111111110011000000000000101101111111111111110000000000000001011111111111101001111111111111001000000000000000000000000000110000000000000010100111111111110110111111111111110001111111111110100000000000000011011111111111111010000000000010111000000000000000011111111111110101111111111101110111111111110001111111111111001101111111111100000000000000000001000000000000010011111111111100011111111111111100100000000001100111111111111111101111111111110111111111111111100100000000000001111111111111100011000000000000011010000000000100000000000000000100100000000000011111111111111101000111111111111010100000000000010110000000000010011111111111111011000000000001101101111111111110110111111111111101111111111111110101111111111110000000000000000000100000000000101011111111111100110000000000000010000000000000101001111111111111001000000000001000011111111111110100000000000000000000000000000000011111111111101010000000000010010111111111110110111111111111100111111111111110110111111111111010100000000000000110000000000010010111111111111001011111111111111011111111111011101000000000000000100000000001010101111111111111000000000000001001111111111111111111111111111111100111111111110100000000000000001111111111111100010111111111110011011111111111101111111111111110100000000000000011000000000000011011111111111101000000000000001000100000000000100101111111111110010000000000000100111111111111100000000000000010011000000000000010000000000000000011111111111011000111111111111111111111111111100011111111111110011111111111111001100000000000000010000000000001100111111111110100100000000000010000000000000010001111111111110111111111111111101010000000000110000111111111111011000000000001000000000000000100101000000000001110000000000000100011111111111111111000000000001001011111111110111100000000000000110111111111111110000000000000000110000000000010111000000000001001100000000000100110000000000010110111111111110010100000000000000111111111111101100000000000000100000000000000101001111111111110011111111111110001111111111111111001111111111111100111111111110000111111111111100000000000000101001111111111111011111111111110110110000000000000101000000000001100000000000000110011111111111100111000000000001101100000000001000010000000000000100111111111110010100000000000100010000000000000101000000000000001100000000000001100000000000011111000000000000000000000000001010010000000000000100000000000000010100000000000010111111111111111101000000000000000011111111111111101111111111110000000000000001000111111111111011011111111111100001000000000000100000000000000001000000000000000010111111111101100000000000000000101111111111110110000000000000000000000000000001110000000000000101111111111111101111111111111011111111111111110111000000000001011011111111111011001111111111110101000000000010000100000000000000101111111111101100111111111111110100000000000110010000000000000010000000000000001000000000000100000000000000000100000000000000100100000000000010001111111111110100111111111111000000000000001000001111111111110011000000000000010111111111111111101111111111101100000000000000001111111111111101100000000000000010000000000000010111111111111100111111111111110111111111111111101011111111111110101111111111110110000000000000101011111111111001110000000000001010111111111110100111111111111011110000000000001001000000000010000000000000000101100000000000100101000000000001011100000000001001110000000000100110111111111110110011111111111111011111111111111001111111111111010100000000000010111111111111111000111111111110001000000000000101001111111111111000000000000000101111111111111100001111111111101110000000000001101000000000000100100000000000001000111111111111110000000000000000111111111111111110000000000000011011111111111001110000000000001100111111111110010100000000000001001111111111101001000000000000110000000000000001110000000000000100000000000001000011111111111111110000000000000010111111111101110011111111110110011111111111101011111111111110001111111111111010000000000000011100111111111111101000000000000011100000000000011000000000000000010011111111111000011111111111111000111111111111010100000000000011010000000000000101000000000001101100000000001001000000000000100100000000000000001100000000000001111111111111110001000000000010011111111111111001111111111111111001000000000000101100000000000000001111111111101111000000000001011100000000000011100000000000000010000000000000101100000000000011111111111111101000000000000000010000000000000010011111111111110100000000000001111011111111111111100000000000100100000000000001010000000000000110000000000000011101000000000100001100000000000101100000000000000111111111111110111000000000000000101111111111101111111111111101011100000000000101111111111111111011111111111111010111111111111101001111111111100100000000000010101100000000000011000000000000001101000000000011001000000000000011010000000000101011000000000001100000000000000101011111111111111000000000000100000100000000001001000000000000011100000000000011101100000000001101100000000000100001000000000011010000000000001011010000000000101110111111111110110100000000000000010000000000000101000000000001010000000000000110101111111111111101000000000001000011111111110110011111111111110001111111111101110000000000000000101111111111110111000000000001100000000000000101001111111111100011111111111111011000000000000010111111111111101100000000000001010000000000000010110000000000010000111111111111010100000000000001000000000000011111111111111111001100000000000010010000000000001111111111111111101111111111111111011111111111101100000000000001011100000000000100110000000000100010111111111111011111111111111100100000000000100000000000000101010000000000011101000000000001100010000000000011011100000000011011110000000001110101000000000000010100000000000100111111111111111110000000000001110000000000011000010000000001001111000000000011001100000000001100110000000000000110111111111111110011111111111110111111111111001110000000000000011111111111111111100000000000010011000000000000110000000000001010100000000000010101000000000000110100000000000110110000000000011001111111111111010000000000000011100000000000001100111111111111101000000000000011101111111111110000111111111111011111111111111111100000000000001101000000000000101100000000000000011111111111100111000000000010001111111111111101001111111111100001000000000010100000000000000001100000000000011101000000000000110000000000000101010000000000010101000000000010001100000000000110100000000000001001000000000000011100000000000001101111111111000100000000000000110011111111110110011111111111100110000000000010101011111111110110101111111111110011000000000000011100000000001001101111111111111111111111111110110011111111101001001111111110100011111111111110111111111111111001111111111111100001000000000011110100000000000100110000000000010011000000000010111000000000011101000000000001010100000000000000111100000000010000100000000000010110111111111101110011111111111101011111111111011001000000000001110000000000001000001111111111111110000000000001001011111111111111010000000000001100111111111111101011111111111100101111111111110001000000000001110100000000000001100000000000000000000000000001000100000000000011010000000000000010000000000001101011111111111110010000000000000001111111111110000111111111111111010000000000011001111111111111111100000000000010111111111111111111111111111111010000000000000011010000000000000001000000000000001011111111111011111111111111101010111111111110010000000000000010010000000000000001000000000000101100000000000010011111111111101001111111111110110100000000000001101111111111110111111111111111100011111111111101111111111111111111000000000000011011111111110111011111111111111011000000000000000000000000000000001111111111110111000000000000100011111111111010111111111111110100111111111111010011111111111101100000000000001101000000000000001100000000000000100000000000010010111111111111000111111111111011001111111111111110000000000000010011111111111101000000000000010001000000000000001111111111111101111111111111111000000000000000101100000000000000001111111111111100000000000000001011111111110111011111111111111111000000000000110111111111111111011111111111111100111111111111011100000000000100101111111111111100000000000010000000000000000000100000000000011110111111111111011011111111111110100000000000001111111111111101101011111111111100100000000000000000000000000000100100000000000000010000000000000011111111111111110111111111111110111111111111110011000000000000100111111111111110011111111111101000111111111110100011111111111111110000000000011010000000000010010100000000000000001111111111110101111111111111010111111111111111000000000000011010111111111110101100000000000000001111111111111101000000000001100000000000000101011111111111111111000000000001010011111111111110101111111111111010111111111111101111111111111110110000000000001110000000000001000111111111111010011111111111100100111111111111010000000000000000101111111111111111000000000000000000000000000101000000000000000101000000000000010011111111111101110000000000001101000000000000000000000000000011001111111111101011000000000000111000000000000010100000000000001001111111111110111000000000000011100000000000001011111111111111110111111111111110000000000000010001000000000001111011111111111100110000000000010101111111111110100111111111111111101111111111101101000000000001000100000000000011101111111111111001111111111110101111111111111101011111111111101100000000000000010000000000000110011111111111101110111111111111010011111111111101101111111111110011000000000000000000000000000100110000000000000100000000000000110111111111111011010000000000010100111111111111000100000000000000010000000000001010111111111111011100000000000111111111111111111000000000000000111011111111111001001111111111101101111111111101111100000000000111001111111111100101000000000000010111111111111101011111111111011110000000000000111100000000000010001111111111111101111111111111010111111111111101001111111111010101000000000001001000000000000000000000000000000101111111111110111111111111111101010000000000000100111111111110100111111111111100000000000000001011000000000000110111111111111111001111111111110011111111111111100011111111111100110000000000001000000000000000000000000000000011011111111111111101000000000000010011111111111101110000000000000101111111111111100111111111111010110000000000000000000000000001000111111111111001010000000000000000111111111111001111111111111100000000000000000111111111111111101100000000000011110000000000000101111111111101111000000000000110111111111111100011111111111101101000000000000000001111111111110101000000000000011111111111111110110000000000000100111111111110111100000000000010001111111111110111111111111111100111111111111010010000000000000001;
endcase
end
endmodule



module lut_weights_4(sbyte,addr);
input [3:0] addr;
output reg [41471:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0100: sbyte = 41472'b000000000000000100000000000010000000000000101111000000000000000000000000000110000000000000010100111111111111001111111111111000011111111111110010000000000000100100000000000000001111111111110001000000000000000000000000000011000000000000010001111111111111110011111111111111010000000000000011000000000000000011111111111100100000000000000110000000000000011111111111111100011111111111100111111111111111110111111111111100000000000000000000111111111111100111111111110110110000000000000000111111111110010000000000000100000000000000010010000000000000000000000000000100100000000000001110111111111111011000000000000000001111111111111001111111111110111000000000000001001111111111101011000000000000001100000000000011011111111111011100111111111110101111111111111010000000000000010110000000000000010011111111111110000000000000010011111111111111011100000000000010000000000000000110000000000000001100000000000001000000000000000101000000000001011111111111111101011111111111111101000000000000000000000000000001000000000000001010111111111110111011111111111111001111111111111100111111111101111000000000000010110000000000110000111111111110110000000000000110010000000000000111000000000010110011111111111110010000000000000110000000000001111000000000000011111111111111110001000000000011100000000000000000001111111111111111111111111110011011111111100001101111111111001101111111111100010011111111111001000000000000110100111111111101101000000000000111110000000000101000000000000001011100000000000101001111111111101110111111111111110011111111111100111111111111111110111111111111011100000000000001010000000000001000111111111110011100000000000010001111111111110010000000000000100111111111111110101111111111111100000000000000011011111111111110110000000000001110000000000000000000000000001000111111111111011111000000000010010111111111111110001111111111011111000000000000010011111111111111111111111111101010111111111111100011111111110111110000000000110000111111111111001100000000000100010000000000011111000000000010010100000000000111011111111111111010000000000000101100000000000001111111111111101100111111111111010111111111111010110000000000001101111111111110111111111111111100011111111111111000000000000000000011111111111110100000000000001100111111111111010100000000000110100000000000000001111111111111111100000000000000100000000000011010000000000000000000000000000000101111111111111100000000000001000100000000000000110000000000001101111111111111000100000000000010011111111111111010000000000000010000000000000010010000000000000111000000000000111111111111111100011111111111100111111111111101101100000000000000001111111111101001000000000000111000000000000001101111111111011011111111111110110100000000000100000000000000000100000000000000011000000000000011101111111111111011000000000000101000000000000001000000000000000010000000000000011100000000000010110000000000000010000000000000001011111111111101011111111111110100000000000000100000000000001000111111111111111101000000000010010100000000000101111111111111100111000000000000001011111111111111001111111111110010111111111110010111111111111101100000000010000100000000000000000000000000000110101111111111010010111111111111101011111111111011111111111111110010000000000010000100000000000010000000000000000001000000000001010111111111111111000000000000000000111111111111111000000000000000000000000000010001111111111110100111111111111111101111111111111001111111111111000000000000000000101111111111110101000000000000001000000000000011110000000000001111000000000001000100000000000011100000000000011101111111111111101000000000000100001111111111101111000000000001010100000000000110001111111111111111111111111111101100000000000011000000000000100001111111111111100111111111111101001111111111111011111111111110110111111111111100101111111111111110000000000000111011111111111110100000000000001111111111111111011111111111111100111111111111111110111111111111011111111111111011111111111111110000111111111110110011111111111111100000000000001111111111111110101000000000000101010000000000000011000000000000100011111111110111101111111111110110111111111111101100000000000010011111111111111001111111111110000100000000001001000000000000000001111111111111001000000000000000010000000000000100000000000001001000000000000100100000000000010111111111111111000011111111111110011111111111100101111111111111001100000000000010001111111111100110111111111111011100000000000001100000000000000000111111111111101100000000000000101111111111110101000000000000001111111111111111001111111111111011000000000000001011111111111101110000000000000001111111111100111000000000000000001111111111111011111111111110110111111111111100111111111111111001000000000011010000000000001001100000000000100000000000000010111000000000001000000000000000011011000000000001010100000000000011101111111111111010000000000000111000000000001010010000000000000011111111111110100000000000000010111111111111111110111111111101111111111111101100111111111110010100111111111111011111111111111100000000000000000011000000000000111111111111111010111111111111111101111111111111100011111111111110001111111111111101000000000000000011111111111110011111111111110100000000000000000011111111111101110000000000000100111111111111100100000000000010010000000000000010000000000001000000000000000000000000000000001000111111111110010111111111111100110000000000000100000000000010000100000000000100100000000000001011111111111110100100000000000011101111111111110000000000000001000011111111111101011111111111011011000000000000111000000000000000000000000000000101000000000000000111111111111001000000000000011000000000000001010000000000000100001111111111111010000000000000001100000000000010011111111111101100000000000000101100000000000011111111111111110010000000000001101111111111111000010000000000010010111111111110011111111111111100110000000000001011000000000001000011111111111100001111111111111100000000000000000100000000000000101111111111101010111111111111110111111111111001011111111111110111000000000001101100000000000000111111111111111011000000000000010100000000000011000000000000001111111111111111110011111111111011111111111111111111000000000000011100000000000000101111111111110000111111111110111100000000000001100000000000011111111111111111110000000000000001101111111111111001111111111111101111111111111011101111111111101011000000000000101100000000000101101111111111111110000000000000000111111111111011110000000000011100000000000000110111111111111100100000000000010100000000000000011000000000000000000000000000001101000000000001010100000000000011011111111111101000111111111111010111111111111011011111111111101110000000000001110111111111111010000000000001001011111111111101001111111111111001010000000000010001000000000000111111111111111011011111111111110010000000000000010111111111111011001111111111110001000000000000100111111111111100111111111111110010000000000001101100000000000001101111111111101110111111111111101011111111111101111111111111111000111111111111010011111111110101110000000000010011111111111111010011111111110101010000000000001100000000000001111000000000001100110000000000010010000000000000110011111111111111000000000000010011111111111111101100000000000100101111111111110100111111111101111100000000000011111111111111110010111111111110100111111111111101111111111111111010111111111111110100000000000010100000000000000010111111111111010100000000000001001111111111110101000000000000100100000000000010001111111111111011000000000000001011111111111111001111111111100011000000000000011100000000000001111111111111110010000000000001110100000000000001011111111111111100111111111111001100000000000001100000000000000011000000000001011111111111111101001111111111110011000000000000000100000000000010000000000000001011000000000000101000000000000000011111111111110111000000000001111011111111111100011111111111111011000000000001010011111111111111011111111111111111111111111111011011111111111100000000000000011000000000000000011011111111110111001111111111111110000000000000111011111111111111110000000000010000000000000000010111111111111111111111111111111110000000000000111011111111111011110000000000000101000000000010010111111111111111001111111111110000111111111110100000000000000010100000000000010010111111111101111111111111111010010000000000100000111111111110000000000000000000000000000000000011000000000000110111111111110010011111111111011111000000000010011111111111111000001111111111111111000000000101110000000000001100001111111111101001111111111111110000000000000010111111111111111110111111111111011100000000000101001111111111100011000000000001000111111111111111101111111111111110111111111110111111111111111001010000000000000100000000000000001000000000000010001111111111111111111111111111010100000000000100101111111111111100111111111111001111111111111000101111111111111001111111111111011100000000001010100000000000100110000000000001101000000000000100101111111111110110000000000000110000000000000111001111111111110100111111111111100111111111111001100000000000010111000000000000000000000000000000000000000000010110000000000000111111111111111101111111111111111000000000000001010111111111111111011111111111111001111111111111001000000000000000000000000000010110000000000001010000000000000001011111111111110011111111111110000011111111111101100000000000001000111111111111111000000000000101100000000000010110000000000001000111111111111011010000000000001000111111111111110100000000000100100000000000001100000000000000001111111111111011100000000000011111111111111111101011111111111011101111111111101101111111111110100000000000000000111111111111111010000000000001101100000000000100001111111111100000111111111110101111111111111110001111111111111101000000000000011100000000000010000000000000000110111111111111110111111111110100111111111111101101111111111111010011111111111100101111111111110110111111111110011011111111111110011111111111111011000000000001000100000000000010110000000000000110000000000000011000000000000010000000000000010100000000000001000000000000001000111111111111110111000000000001011000000000000001111111111111111011111111111110110011111111111100101111111111101010111111111011111011111111110101011111111111110011111111111101110100000000010000010000000000000101000000000001101100000000000010100000000000000000111111111111110100000000000001011111111111111001111111111110110100000000000000010000000000000001111111111111001111111111111101010000000000001001000000000000101100000000000010010000000000011010000000000000101000000000000011011111111111111001111111111111011011111111111101100000000000010010111111111110010100000000000100110000000000011100000000000001110000000000001011101111111111101000000000000000011100000000000000101111111111101010000000000010100100000000000001000000000000001111111111111111101000000000000001110000000000000110111111111111110000000000000001000000000000001000000000000000010011111111111011110000000000000101111111111111001000000000000000000000000000011010000000000001110111111111111010101111111111011010000000000001001111111111110001010000000000010010111111111110111000000000000001010000000000001110111111111111111111111111111111010000000000000010000000000001110011111111111100011111111111101011000000000000101000000000000000010000000000011110111111111111001111111111111100110000000000010001111111111110010000000000000000100000000000000100000000000000001100000000000001001111111111101110111111111111100111111111111101010000000000011111111111111111101000000000000011010000000000000001000000000000011100000000000001100000000000000001000000000000010011111111110100000000000000100111111111111111111111111111111101001111111111110111111111111110111111111111111101100000000000001001000000000001000100000000001000000000000000100001000000000001010000000000000111010000000000000111000000000001110000000000000100101111111111111011000000000010011111111111101100001111111111100011111111111110100111111111101111010000000000011110111111111011111000000000000101110000000000100011000000000000000100000000000000010000000000001111000000000001000000000000000000110000000000000000000000000001100100000000000000111111111111110100111111111111111100000000000010110000000000010001111111111111111000000000000001100000000000000110111111111111111111111111111110100000000000000010000000000010010000000000000101111111111111100000111111111110101111111111111001001111111111111010111111111111100011111111111011111111111111011101000000000000100000000000000000110000000000101010000000000000010000000000000101001111111111110110111111111111110111111111111111111111111111110011000000000000000111111111111111001111111111111011000000000000001100000000000000111111111111111110000000000000010100000000000001001111111111111100000000000000100100000000001000000000000000010100000000000001100011111111111011001111111111101010111111111100001011111111111100101111111111100100000000000000101111111111111101011111111111111011000000000000111111111111111001110000000000001001111111111111111100000000000011010000000000000101000000000000010011111111111101000000000000001001000000000000000111111111111100101111111111100010111111111111001011111111111110001111111111110011000000000000101011111111111101010000000000000000111111111110111011111111111001000000000000001101000000000000001100000000000000111111111111110000111111111111011100000000000010011111111111101011000000000000110011111111111111010000000000000000111111111111011000000000000000001111111111111000111111111111101111111111111000011111111111100100000000000001111000000000000100100000000000010011000000000011001000000000000110010000000000101000000000000100111000000000001011100000000000010111000000000011111011111111111111111111111110110110111111111100000011111111110011001111111111010100000000000000100000000000000100010000000000001011111111111111011011111111111011111111111111110101111111111111110011111111111100100000000000000011111111111111111000000000000100111111111111111010111111111111100011111111111111110000000000000000000000000000001111111111111001110000000000001100111111111110111100000000000000011111111111111010111111111111100111111111111110010000000000000100111111111111011111111111111111011111111111111110000000000001011100000000000000001111111111111101111111111111111011111111111100100000000000001010111111111111101011111111111111000000000000000110111111111111011011111111111100110000000000001011111111111111111111111111111111111111111111111100000000000000101011111111111100110000000000001000000000000000001100000000000001000000000000001010111111111111111100000000000011000000000000001001111111111111110111111111111011110000000000001100000000000001110111111111111101001111111111110101111111111111111000000000000100101111111111111100000000000001001100000000000000101111111111111011111111111111101100000000000010011111111111111010000000000000011100000000000000000000000000000111000000000000000111111111111011111111111111111111111111111110011000000000000110010000000000010111111111111111001000000000000000110000000000000001111111111111100111111111111010000000000000001001111111111111110000000000000001111111111111111001111111111110110100000000000000001111111111100111000000000000010111111111111110110000000000000000111111111111111111111111111101110000000000000000111111111111010000000000000010100000000000010011000000000000001100000000000000010000000000000001111111111111100011111111111101010000000000011011111111111111110100000000000011101111111111101011111111111111011011111111111010111111111111111001111111111111111100000000000111011111111111111101000000000000110011111111111101011111111111111100111111111111000111111111111011011111111111110101000000000000001100000000000101000000000000011100000000000001000000000000000010100000000000000000111111111111111000000000000000101111111111110111000000000001010100000000001001101111111111100001000000000001001000000000000101110000000000001001111111111111100000000000000000000000000000001000000000000000001011111111111100101111111111101100111111111111010111111111111111100000000000000010000000000001000100000000000001011111111111111000000000000000011000000000000000101111111111111110000000000001011111111111111010110000000000000000111111111111000100000000000000001111111111110100111111111111100111111111111101011111111111110010000000000000111000000000001000011111111111111010000000000001111111111111111001111111111111110010111111111111011111111111111010011111111111101101000000000001010111111111111100001111111111110100000000000000101100000000000001110000000000000011000000000000111011111111111110001111111111011010000000000001011000000000000010101111111111101110111111111111111111111111111101111111111111111000111111111110101011111111111011011111111111101011000000000000000000000000000101101111111111110101000000000000011011111111111100000000000000000101111111111101001111111111111010011111111111010001000000000001000000000000000100101111111111100000000000000000110100000000000001000000000000000000000000000011111100000000001000100000000000000000000000000011000100000000001011010000000000000001000000000011000100000000000101110000000000000000111111111011101111111111110000011111111110001011000000000100001000000000010000111111111110111100000000000001111000000000000110001111111111010110111111111111001100000000000000101111111111110001000000000001001100000000000011011111111111111001111111111111101011111111111111101111111111111010000000000001011011111111111111101111111111110101000000000000000000000000000011011111111111100101000000000000100111111111111111011111111111101100000000000000101100000000000111101111111111110110000000000000011100000000001110010000000000011011111111111111111011111111111100011111111111101010000000000001001100000000000000010000000000000001111111111111001111111111111011100000000000010100111111111111110011111111111101001111111111111100111111111111110000000000000101010000000000000101000000000001101000000000000010010000000000001110000000000000110000000000000001010000000000010101111111111111101000000000000011011111111111111101000000000000001100000000000100110000000000000000000000000000100100000000000011111111111111111010000000000000010011111111111101111111111111111001000000000001011100000000000101000000000000001010000000000001000111111111111111000000000000010101000000000000001011111111111101010000000000001010111111111111100000000000000100111111111111111001000000000001010111111111111101011111111111101010111111111111010011111111111111101111111111111111000000000001000000000000000100001111111111111001000000000000010111111111111100010000000000001000000000000000110011111111111111011111111111010110000000000000000100000000000001100000000000001100000000000001010100000000000100011111111111110110000000000000111011111111111010100000000000001101111111111111011011111111111110000000000000001000000000000000110111111111111011011111111111110010111111111110110111111111110101101111111111100100000000000001001100000000000010011111111111011101000000000011011000000000001001100000000000001110000000000001100000000000000011000000000000000010000000000000011011111111111101111111111111100100000000000000010011111111111110110000000000001011111111111111010011111111111101110000000000000011000000000000100011111111111110100000000000000011000000000000000000000000000000000000000000000001000000000010111011111111110101100000000000001010111111111111010011111111111101001111111111111000000000000001001011111111111111110000000000011111000000000010000111111111111111001111111111100001000000000000111111111111111111111111111111101101111111111111110100000000000010011111111111111100000000000000011100000000000000110000000000000011000000000001010111111111111111011111111111111001111111111111011000000000000101101111111111110110000000000001001000000000000001111111111111010000000000000001000011111111111110101111111111010111000000000010000000000000000000001111111111110111000000000000001011111111111011010000000000000011000000000000001100000000000001011111111111111000000000000000001100000000000010100000000000000000000000000001000100000000000000000000000000000110000000000001001011111111111010011111111111110010000000000000001100000000000000001111111111110011111111111111010100000000000001100000000000010001000000000000110100000000000010010000000000000010111111111111110100000000000011001111111111110011000000000000011111111111111101001111111111011100000000000010000111111111111001101111111111110000000000000000001100000000000001011111111111110100000000000000100100000000000000100000000000110010111111111111110000000000000011100000000000011011000000000000011000000000000110010000000000001010000000000011101011111111101011001111111101111100000000000011010011111111101101011111111110101000000000000101000000000000000011001111111111010010111111111111010111111111111110110000000000010001111111111111010111111111111101001111111111110111111111111110001100000000000000000000000000000100000000000010100000000000000011110000000000000000000000000000100111111111111111111111111111111100000000000001000011111111111111110000000000000111000000000000111000000000000011101111111111111100000000000001001000000000001000100000000000000000000000000010100000000000000010010000000000001110000000000001001100000000000000011111111111111001000000000000010011111111111101001111111111100001000000000000101011111111111110101111111111110010111111111110101111111111111111011111111111111001000000000000010100000000000001101111111111111111000000000001010011111111111010000000000000000011000000000001010011111111111100001111111111101111000000000000000000000000000100011111111111110101000000000000111000000000000110001111111111010101111111111111001111111111111011101111111111101100000000000000100000000000000001101111111111110111000000000000000111111111111110010000000000000101111111111111001011111111110100000000000000000100000000000000100000000000000010001111111111110001111111111111100011111111111011011111111111111110000000000000101000000000000000001111111111011111000000000001001000000000000000001111111111101111000000000000101111111111111111000000000000000111000000000000010011111111111000101111111111100111111111111111011100000000000010001111111111101001000000000001011100000000000101011111111111100111000000000001011100000000001011000000000000011001000000000000101000000000000011110000000000011000000000000000101100000000000001101111111111110101111111111111101111111111101110011111111110111001111111111110011111111111110111111111111111000010000000000100111000000000000111111111111111001010000000000001011000000000000001011111111111111100111111111110000111111111111011010000000000000110000000000000000111111111111111100000000000001000000000000000010011111111111110101111111111111011000000000000001100000000000001100000000000001011111111111110011000000000000001010000000000000001000000000000010011111111111101100000000000000011111111111110011011111111111011000000000000000111000000000000010000000000000111010000000000010101000000000001010100000000000100101111111111111001111111111111001011111111111100010000000000000000111111111111010011111111111101001111111111110111000000000000000111111111111101101111111111111110000000000000000011111111111100111111111111110011000000000000010100000000000001101111111111111111111111111111100000000000000001101111111111100010000000000001010000000000000011001111111111100111000000000001110000000000001001000000000000000000111111111111110011111111111110101111111111111101000000000001000000000000000011100000000000000100000000000000011000000000000001101111111111110011000000000000101011111111111011010000000000000000000000000001000100000000000001111111111111111010000000000001100111111111111111011111111111101110000000000001001011111111111000011111111111111011000000000000101011111111111001101111111111111000000000000000011111111111111111111111111111101110000000000000000011111111111101101111111111100110000000000000111000000000000010111111111111101011000000000000100100000000001000101111111111111101111111111110111000000000000001001111111111111111111111111111100011111111111110000000000000010111111111111111011011111111111011100000000000000110111111111111110011111111110101101111111111010100000000000100100000000000000010001111111110111111000000000000111000000000001100000000000000001011111111111111111000000000000001100000000000001111111111111111101011111111111111100000000000001011000000000000001000000000000000010000000000000100111111111111110000000000001001011111111111110110111111111111001011111111111010101111111111101111111111111111101111111111111111011111111111110001111111111111100011111111110011111111111111010010000000000001001000000000000000000000000000000010111111111111101100000000000101010000000000011101111111111101101000000000000000011111111111101101000000000000100011111111111001011111111111110101000000000000001100000000000010100000000000000001000000000001101111111111111110110000000000001110000000000000010100000000000001100000000000000111000000000000110000000000000000101111111111111010111111111110101100000000000111001111111111110111111111111111110011111111111111001111111111100010111111111111100011111111111110100000000000011001000000000000000000000000000100011111111111101111111111111111110100000000000010111111111111111111000000000000100011111111111101101111111111110010111111111110100011111111111111011111111111110111000000000001100011111111110111101111111111110101000000000000001100000000000110010000000000000011111111111111110111111111111101101111111111111001000000000000111111111111111111100000000000000101111111111111110111111111111100001111111111101100111111111111110011111111111100001111111111111110111111111111011011111111110110011111111111110000111111111111101000000000000011100000000000010000000000000000000011111111111100001111111111111100000000000001010100000000000001010000000000010001000000000001010111111111111110001111111111111010111111111111110000000000001101100000000000000001111111111110100111111111101000101111111110100111000000000000011100000000010000000000000001001111000000000000001111111111111111001111111111101010111111111111111100000000000000011111111111111000000000000000001100000000000000001111111111110111000000000000110000000000000010000000000000000001000000000000000011111111111100011111111111101011000000000000010111111111111011010000000000010001111111111111111111111111111101110000000000000110000000000000011111111111111101011111111111100001111111111111110111111111111101000000000000001110111111111111010000000000000001100000000000001101111111111110010111111111111100001111111111111101111111111111101111111111111100010000000000000000000000000001001011111111111101101111111111111100000000000000101011111111111101010000000000001010111111111111101100000000000100000000000000000001000000000001000100000000000000110000000000100101111111111111100011111111111011011111111111010011111111111111010111111111110111001111111111101100111111111111111111111111111101000000000000010010111111111111011011111111111110000000000000000110000000000001100100000000000001011111111111110011000000000000010111111111111110011111111111110011111111111110010011111111111001111111111111100011111111111111001100000000000100001111111111111000000000000000111011111111111010100000000000010000000000000001000111111111111011010000000000001101111111111111101111111111111111111111111111110100000000000001010000000000000011000000000000000000111111111111011011111111111010010000000000000111111111111111111011111111111111010000000000001001000000000001011111111111111111111111111111111110000000000011011111111111111110100000000000001100000000000001011111111111111101000000000000000000000000000000110100000000010101000000000000110001111111111011011011111111111010111111111111110101111111111101011111111111110101111111111110111000111111111111111011111111111111100000000000000000111111111101100100000000000001010000000000001100111111111111010000000000000000001111111111100111000000000000011000000000000000000000000000001100111111111111111011111111111111001111111111111101000000000000001111111111111111110000000000001010000000000000011100000000000000110000000000000111111111111111011000000000001000100000000000100011111111111110001111111111110001101111111111101111111111111111010111111111111001011111111111100010000000000000000111111111111010111111111111110000111111111111101111111111111110101111111111100111000000000000000011111111111111000000000000000001000000000000011011111111111100011111111111111101000000000000011111111111111010010000000000001100000000000000111111111111111100011111111111110001000000000000011100000000000001101111111111111010111111111111011011111111111111000000000000000101000000000000000000000000000001010000000000011001000000000000111011111111111111000000000000001001111111111111111011111111111111001111111111110000000000000010000111111111111100000000000000010011000000000000000000000000000001001111111111111010111111111111100111111111111100000000000000001010111111111111001111111111111010110000000000000011111111111111010011111111111100111111111111100000000000000001001100000000000011010000000000100100000000000000101111111111111101101111111111011000000000000000000000000000000111100000000000010001111111111111000100000000000011010000000000001111111111111110000011111111111100110000000000001000111111111111111011111111111010110000000000010000111111111111110111111111111001111111111111111011111111111111100111111111110011001111111111001110000000000010111000000000001011000000000000110100111111111101000000000000001001000000000001011111000000000000000100000000000011000000000000001110000000000000011011111111111001011111111111111011111111111111101000000000000010101111111111101101000000000001011011111111111111000000000000011000111111111110011011111111111101111111111111100111000000000000000011111111111101001111111111101110000000000010100111111111110100101111111111011100000000000000111100000000000110110000000000101001111111111110001111111111111100010000000000100100111111111110001111111111111110000000000000000000000000000000100100000000000001100000000000000000111111111111101111111111111011011111111111110000111111111111111100000000000000001111111111111111111111111111011100000000000001101111111111110000000000000001101111111111111111110000000000000100111111111110111011111111111001111111111111011101000000000000110100000000000011110000000000001001111111111111111000000000000000000000000000001100111111111111111011111111111101100000000000010101000000000000011000000000000001011111111111011010111111111110110100000000000000111111111111111011111111111111001111111111111001011111111111100010111111111111101100000000000000010000000000000000111111111110011111111111111000110000000000001111111111111111111000000000000011100000000000010001000000000000110111111111111101101111111111011010000000000000001100000000000010010000000000000001111111111111100111111111110110111111111111100111000000000000110000000000000000001111111111101000111111111111010100000000000010000000000000010101000000000010110111111111111010010000000000001101000000000011011000000000000011100000000000011010000000000001001011111111111100111111111111101001111111111001110111111111100110001111111110001101000000000001000100000000001000101111111111110010111111111111111100000000010011110000000000111001000000000001100011111111111101110000000000000101111111111111101000000000000001111111111111111010000000000000000011111111111011110000000000010010111111111111100100000000000010100000000000000000111111111111010100000000000000111111111111110110000000000001000111111111111111110000000000000000000000000000000011111111111110101111111111110001000000000000000011111111111100100000000000001001000000000001110100000000000010101111111111111000000000000001000011111111111111001111111111111000000000000001010011111111111011110000000000010110000000000000101111111111110100010000000000000101000000000001001011111111111100101111111111011101000000000001001000000000000000011111111111111010000000000001001011111111111100000000000000001110000000000000000011111111111111100000000000001011000000000000110011111111111110010000000000010001000000000000000011111111111101001111111111111100111111111111011100000000000000011111111111111100000000000000011000000000000011000000000000000101000000000001011011111111111100000000000000000000000000000000001100000000000011110000000000001101000000000000011111111111111001001111111111111011111111111111011100000000000010001111111111110011111111111111110100000000001000110000000000001011000000000000000011111111111101111111111111111100111111111111110111111111111111101111111111101110111111111111111111111111110111000000000000000110111111111111111011111111111111110000000000100001000000000001001011111111110101100000000000000111000000000000111100000000000111001111111111110100000000000000010100000000000111101111111111111111111111111111001011111111111101001111111111110100111111111100000011111111110111010000000001100101111111111101110111111111111011010000000000011001111111111110010011111111111011100000000000100011111111111110111000000000000001100000000000000101000000000000010011111111111111000000000000000011000000000000110111111111111101011111111111110100111111111111010100000000000010110000000000010000000000000000001100000000000001001111111111110000111111111111100100000000000010001111111111111110000000000000111011111111111100111111111111101100000000000001110000000000000111010000000000010100000000000000101011111111111110111111111111110111111111111110100100000000000011101111111111111111000000000000000011111111111111000000000000000000111111111111101100000000001000100000000000010101111111111111011011111111111111101111111111111011000000000000000011111111111110101111111111110110111111111111101111111111111111101111111111111010111111111101110111111111111100111111111111111001111111111110100011111111111111011111111111111000000000000000000100000000000001101111111111110011000000000000110111111111111110011111111111111011000000000000100011111111111101101111111111111101000000000001001011111111111110001111111111111111000000000000100111111111110111101111111111110101000000000000011000000000000011110000000000000001000000000000000000000000000100010000000000011000000000000000000100000000000010011111111111111010000000000000000000000000000010000000000000000111111111111111100100000000000000000000000000010011000000000000000011111111111010011111111111011000000000000000100111111111111101001111111111110000111111111111110100000000000001110000000000000101000000000001100000000000000011010000000000001001000000000011100100000000000100001111111111111001000000000011000000000000000001101111111111101110111111111111011011111111111011010000000000001000111111111111001111111111110101111111111111000101111111111110111000000000001001111111111111111101111111111111110111111111111010011111111111111101000000000000010000000000000001100000000000001000000000000000010011111111111111110000000000000000000000000000011100000000000101000000000000010010111111111111011000000000000010010000000000010110000000000000110011111111111101000000000000001000111111111111001000000000000001111111111111001001111111111110101111111111111101000000000000010111111111111111111000000000000000010000000000100000000000000000000011111111111100110000000000000100111111111110101011111111111101011111111111100111000000000000110000000000000010101111111111101010111111111111011100000000000011100000000000000010000000000000001100000000000000011111111111111100000000000000100111111111111100001111111111110110111111111111001100000000001000001111111111111110111111111110110111111111111101011111111111100111000000000000001100000000000100110000000000011011000000000001000100000000000011101111111111101010111111111111111011111111111100010000000000000001111111111111110111111111111110010000000000010011000000000000000000000000000010111111111111110100000000000000001000000000000100110000000000000000111111111111001011111111111111110000000000010100111111111111101011111111111011100000000000000000000000000000011100000000000110000000000000000101000000000000100100000000000011000000000000010111000000000000001000000000000101001111111111101100000000000000000011111111111110011111111111111110111111111111101100000000000101110000000000011101000000000000010111111111111111001111111111110111000000000000000111111111111110000000000000000111111111111111011000000000000000100000000000000101000000000011000000000000010011011111111111111000111111111101100111111111111101111111111111001101111111111110111011111111111111000000000001000101000000000000010011111111111110110000000000100010000000000001011111111111111111111111111111111000000000000000001111111111111100001111111111101111000000000000100111111111111110110000000000000111111111111110111000000000000000100000000000011011111111111110110011111111111101110000000000000101000000000000011111111111111001111111111111101110111111111111000011111111110111111111111111110001000000000000000000000000000001010000000000000000000000000001000100000000000000110000000000100111000000000000101000000000000110111111111111100111111111111111011000000000000001110000000000001001000000000000111111111111111110110000000000000110111111111110111000000000000000101111111111110101000000000000000011111111111101100000000000001011111111111111110000000000000100011111111111110011000000000001111100000000000011011111111111101000111111111110001111111111111100101111111111111111111111111110101111111111111110010000000000001100111111111111101011111111111101110000000000000011000000000000110000000000000001001111111111111100000000000000001100000000000001001111111111100011000000000001100000000000000000001111111111111000000000000000111100000000000100010000000000001010111111111111101111111111111111110000000000000000000000000000001100000000000100111111111111111000000000000000001000000000000010010000000000000001000000000000100000000000000100001111111111100110000000000010011100000000000101101111111111101111111111111111110011111111111100011111111111111001000000000000101011111111111111110000000000000111111111111110110011111111111101000000000000011001000000000000100000000000000000000000000000000000000000000000100100000000000101111111111110101101000000000101100000000000001010011111111110111100000000000000000000000000000111001111111111100001000000000000110111111111111111101111111111010110111111111111101111111111111110000000000000000000111111111111001011111111111111001111111111111100000000000000010000000000000011000000000000000000000000000001000000000000000011011111111111110110111111111111001000000000000001011111111111110010000000000001110100000000001001001111111111111000111111111111000111111111111110011111111111101111111111111111110111111111111010101111111111111001111111111110111011111111111111000000000000110100111111111110101111111111111101010000000000010100000000000000010111111111111111000000000000010110111111111111110011111111111101010000000000001001000000000000110100000000000000111111111111101011111111111110110111111111111100101111111111111101000000000000000011111111111111000000000000101110111111111111111100000000000001100000000000001110111111111111011111111111111010111111111111111111000000000000101000000000000100001111111111110100000000000001010111111111111101101111111111111010111111111111101011111111111110000000000000011101000000000000101100000000000010101111111111110100000000000000010000000000000001110000000000010000111111111111111100000000000100010000000000000100000000000000011100000000000001110000000000000000000000000000000100000000000001110000000000000101111111111111110100000000000001000000000000010111000000000000011111111111111110100000000000001110111111111110111100000000000001100000000000011111111111111101111111111111111000000000000000010010000000000001010100000000000000101111111111111000000000000001101011111111111011011111111111101101000000000001111011111111111101011111111111110001111111111100111011111111111000100000000001011001111111111101110100000000001110000000000000110010111111111011001011111111110110011111111111111000000000000000011000000000000000011111111111110011111111111111111100000000000000000000000000100010000000000000000111111111111101001111111111101100111111111110001011111111111010011111111111101001000000000000000000000000000010011111111111110000111111111111010111111111111101110000000000000110000000000001000111111111111101011111111111101110000000000000001111111111111011110000000000000100000000000000000011111111111000110000000000001110111111111111011000000000000010101111111111110110000000000011000000000000000001111111111111110100000000000000101000000000000000111111111111110110000000000000010011111111111101110000000000001010000000000000000000000000000010010000000000000101111111111111001000000000000000111111111111111100000000000001000000000000000010101111111111111110000000000010100011111111111100011111111111111010000000000000111011111111110101111111111111110111111111111111000000000000000011100000000000000000000000000010010000000000001001001111111111110011111111111110011100000000000000000000000000000010111111111111101011111111111100111111111111100000000000000000111111111111111001011111111111111010111111111111100111111111111100110000000000000111111111111111110011111111111101110000000000000011000000000000001000000000000100010000000000001010000000000000001011111111111111001111111111110011000000000000100011111111111111011111111111111011000000000000011011111111111010001111111111011101111111111111010011111111111000011111111111110011000000000001001111111111110110100000000000001111111111111111110000000000000000011111111111111110000000000000010100000000000000000000000000010011000000000001101100000000000000001111111111001011000000000011000011111111110011101111111111010100000000000010010011111111101101101111111111101000000000000000111100000000000001000000000000000111000000000000100111111111111110111111111111111011111111111101110100000000000000000000000000000100111111111111101100000000000110101111111111111110000000000000101100000000000101001111111111111010000000000000001011111111111100011111111111111111;
endcase
end
endmodule



module lut_weights_5(sbyte,addr);
input [3:0] addr;
output reg [82943:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0101: sbyte = 82944'b000000000000111111111111111001101111111111011001000000000010001011111111111011101111111111101010000000000000111111111111111111010000000000000000000000000001101000000000001001110000000000001110000000000001000111111111111001111111111111101100000000000000110111111111111110110000000000000100000000000001010011111111111101010000000000000000000000000000111100000000000010001111111111110000000000000001010111111111111011111111111111011101000000000001011111111111111111111111111111110110000000000000110011111111111111100000000000001000111111111111011111111111111111100000000000011010111111111111100011111111111101010000000000011100111111111101110011111111111111110000000000100011000000000001010111111111111010101111111111111110111111111111110011111111111111011111111111100111000000000000110111111111111111011111111111101010000000000010001111111111111111010000000000001101000000000001000011111111111101001111111111101010000000000011001000000000000000001111111111111001000000000001101000000000000001111111111111111011000000000000010100000000000110010000000000000000000000000000011011111111111100011111111111011001000000000001111011111111111111100000000000010101000000000000011100000000000100101111111111111110000000000000000100000000000001011111111111111101000000000000000011111111111011110000000000000100000000000000000011111111110001001111111110100101000000000000101000000000000000000000000000001111000000000001100111111111111101110000000000001111000000000000101000000000000001000000000000000011111111111111001000000000000010000000000000000100111111111110111011111111111101000000000000010100000000000000000011111111111110011111111111110111000000000001010000000000000111111111111111110000111111111111101011111111110010111111111111100010111111111111001111111111111100001111111111011000000000000001010000000000000111000000000000100110000000000001101011111111111010011111111111111011000000000000000000000000000001101111111111111110111111111110101100000000000101010000000000100000111111111110100111111111111101110000000000001010111111111110100000000000000000100000000000000010000000000000111000000000000010010000000000000010000000000000100011111111111110100000000000000001111111111111111011111111111111010000000000010101000000000000000111111111111000010000000000000100111111111111100000000000000010101111111111110111111111111111010011111111111100000000000000001001111111111110010100000000000001110000000000011000111111111110110111111111111110000000000000010001111111111110100011111111110001011111111110111101000000000000000011111111111101110000000000001100000000000000000111111111111111010000000000000011000000000010000000000000000000000000000000000001000000000000100011111111111100011111111111111100000000000001000100000000000111100000000000000111000000000001010111111111111010101111111111111011111111111111110111111111111110000000000000000000000000000001101111111111111111110000000000000011111111111110001000000000000101010000000000100101111111111110101100000000000101010000000000000110111111111111010011111111111110000000000000001000111111111111011100000000000110000000000000001001000000000000000000000000000101000000000000000000111111111111011100000000000001110000000000010101000000000100010100000000001010000000000000001010000000000000110111111111110111001111111111101001111111111110100100000000000001100000000000000110000000000001011011111111111101011111111111110110111111111111111111111111111110001111111111111111000000000000111111111111111100001111111111111100111111111110110111111111111011000000000000010000111111111111101011111111111100101111111111111100000000000001111000000000000001110000000000000101111111111110001100000000000010000000000000000111111111111110111011111111111101110000000000000011111111111111001100000000000100111111111111111011000000000000000000000000000110011111111111110111111111111111011000000000000100101111111111111101111111111111100100000000000000011111111111110010111111111111111100000000000011011111111111111011111111111110111011111111111101110000000000000010000000000000000011111111111111010000000000000111111111111111101100000000000010100000000000000011111111111111111100000000000000000000000000010100000000000000010011111111111110001111111111110011000000000010010011111111111101011111111111111011000000000000111011111111111110101111111111111011111111111111101000000000000001100000000000000010111111111111111100000000000111110000000000011010111111111111100100000000000001100000000000001111111111111111010011111111111110100000000000001010000000000000100100000000000001000000000000000011000000000000000100000000000000101111111111110110111111111111011000000000000010011111111111111010111111111110110011111111111101001111111111111100000000000000111111111111111110010000000000000000111111111111111011111111111110001111111111110010000000000000100100000000000000001111111111100111111111111111101100000000000000101111111111110010111111111111110100000000000000001111111111110111111111111110111100000000000000101111111111111000000000000000100011111111111111010000000000011000111111111111100100000000000001100000000000010000111111111111101111111111111010011111111111110111000000000000010000000000000001110000000000001000111111111111011111111111111110111111111111110100111111111111101000000000000010010000000000000001000000000000001000000000000010001111111111110010000000000000010011111111111100000000000000010001111111111111101100000000000000010000000000010001000000000001000000000000000000001111111111101010000000000000100000000000000000111111111111111110000000000000100111111111111011100000000000000011000000000000000111111111111110101111111111111011111111111111111011111111111110000000000000001100000000000000000011111111111101011111111111111001111111111111100100000000000010101111111111111111111111111111001000000000000000011111111111111001111111111111110000000000000011011111111111111000111111111111000000000000000000001111111111110100000000000001100111111111111110100000000000001011111111111111110000000000000001011111111111111101111111111110101000000000000000001111111111111100111111111110100100000000000010001111111111111101000000000000011111111111111110001111111111110101000000000000010011111111111111001111111111111011111111111111111011111111111111011111111111101111111111111110110100000000000100011111111111111100111111111110101011111111111111101111111111111111000000000000000111111111111010110000000000000000000000000001000111111111111111100000000000001101000000000000001011111111111101010000000000001010111111111111111000000000000000000000000000000111000000000001001111111111111111100000000000000000000000000000001100000000000101010000000000000101111111111111111111111111111011010000000000001010111111111111110111111111111101000000000000000000111111111111101011111111111111001111111111110010000000000000001011111111111111111111111111110001000000000000110111111111111111110000000000000101000000000000100111111111111100110000000000000000000000000000001011111111111110111111111111111000000000000000011100000000000100000000000000011100000000000000001100000000000011110000000000000111111111111101010111111111110011001111111111100110111111111111011011111111111110101111111111110000111111111111011111111111111110101111111111101100000000000000110000000000000001010000000000000100000000000000001111111111111101110000000000001110000000000000111000000000000100001111111111110010000000000011001000000000001011000000000000011110111111111111010000000000000000011111111111110011000000000001100100000000000101011111111111111000111111111110001011111111111101010000000000000001111111111101100111111111111100010000000000110001111111111101111011111111111111010000000000001100000000000000010100000000000010111111111111100100000000000000010111111111111111000000000000000101111111111110110111111111111011001111111111101101000000000000010100000000000010011111111111111101111111111111100100000000000010100000000000001110000000000000010111111111111111111111111111111011111111111111111111111111111011011111111111110100111111111110111100000000000001100000000000000000111111111111110000000000000000000000000000010000111111111111011011111111111100010000000000100011111111111111011000000000000000001111111111111001111111111110111011111111111110100000000000001010111111111110110000000000000100010000000000000110000000000000110111111111111110011111111111101011000000000001001111111111111100011111111111110011000000000010101000000000000110010000000000001110111111111101110011111111111100000000000000011110111111111100011111111111111111000000000000000101000000000000101111111111111110111111111111101110000000000001000011111111111110000000000000000111111111111111110100000000000010000000000000001110111111111111010111111111111111011111111111100110111111111111111100000000000000001111111111110111000000000001010011111111111010011111111111110100000000000000010000000000000010101111111111111010111111111101001000000000000100010000000000000101000000000000000000000000000101100000000000011000000000000000010111111111110110011111111111110011111111111111001000000000000001000000000000001100000000000000011011111111111111100000000000000001000000000001101111111111111110100000000000010101111111111110111111111111111101001111111111111000000000000000001000000000000001000000000000000001000000000010010000000000001101010000000000101000000000000000110011111111111111111111111111111110111111111101011111111111111100110000000000010001111111111100101111111111110001001111111111111111111111111111011111111111111110101111111111110110111111111110011000000000000010110000000000000110000000000010001011111111111000101111111111111010000000000000001100000000000000001111111111110011000000000000010000000000000101101111111111101000000000000010001011111111111110000000000000001001000000000000100100000000000000010000000000000000111111111111010100000000000001010000000000000111000000000010011100000000000001111111111111111100000000000000011100000000000000001111111111101110111111111101110111111111111011000000000000001001111111111110111111111111110111000000000000010110000000000000010100000000000100010000000000001110111111111110110111111111111111100000000000000101111111111110011011111111101110101111111111101101000000000000001100000000000011100000000000000110000000000001000000000000000101000000000000000101111111111110000011111111111010111111111111101111000000000000000011111111111110111111111111110101111111111111100111111111111101111111111111101111111111111101111011111111111100101111111111110100111111111111100011111111111111101111111111100011111111111110100100000000000000000000000000001001000000000010011100000000001011001111111111111110111111111110111011111111111111100000000000011001111111111111100100000000000011011111111111011000111111111111111111111111111101010000000000011101000000000001101000000000001000001111111111111110000000000001010100000000000000011111111111111100111111111111000111111111111001111111111111101001000000000001010111111111111110101111111111110000000000000000000100000000000000100000000000000001000000000001000011111111111101111111111111011111111111111110110011111111111110000000000000000001000000000000100011111111111010011111111111110001111111111100000111111111110111101111111111011101000000000001000111111111111001001111111111110100111111111111011000000000000101110000000000010100000000000001011100000000000100010000000000011101000000000001001000000000000001000000000000000001111111111111010011111111111111111111111111111001000000000000110100000000000111000000000000010111111111111111001111111111111100010000000000010000111111111111100000000000001011000000000000000011000000000000111000000000001000011111111111111000111111111111010111111111111110111111111111111001000000000000101000000000000000001111111111110101000000000001100100000000000011010000000000000111000000000001100111111111111110000000000000000101000000000000100100000000000011001111111111111000111111111111000011111111111011111111111111100110111111111111010000000000000000011111111111010110000000000000101111111111111100011111111111101100111111111110101100000000000000100000000000001001000000000001010100000000000101010000000000001111000000000000001100000000000001101111111111101010111111111101011111111111111001010000000000000000000000000001000000000000000011111111111111101101111111111111100111111111111111000000000000001001111111111110110011111111111011111111111111101010000000000000100000000000000101111111111111111101000000000000010011111111111011011111111111100101111111111110000111111111110110011111111111100101000000000000100111111111111111010000000000000011000000000010000100000000001010111111111111111110000000000001101000000000000111000000000000001111000000000001100011111111110110101111111111100000000000000010011100000000000000101111111111101000000000000001011100000000000101101111111111101111111111111110111011111111110110111111111111000111111111111110000111111111110111101111111111110110000000000000000100000000000101010000000000000111111111111111100000000000000010101111111111101001000000000001111000000000000101101111111111111000000000000010000000000000000100010000000000001110000000000000101100000000000100110000000000100011000000000000110000000000000010101111111111101100111111111111000111111111110100001111111111011110000000000000000111111111111111011111111111101001000000000011001100000000000001010000000000000001000000000000101011111111111010001111111111111000111111111110010111111111111011100000000000011100000000000000000100000000000110011111111111111101000000000011011000000000001010011111111111100010000000000000101100000000001001010000000000010010111111111111100011111111111101111111111111111001111111111110010011111111111000001111111111011001000000000001101100000000000110010000000000011000000000000010000011111111111000011111111111000110111111111111111011111111110111101111111111110100111111111111011000000000000010110000000000101101111111111111010100000000000000110000000000010000000000000000011000000000000001010000000000001010000000000000100100000000000011000000000000000000000000000000100100000000000000000000000000010100111111111111010000000000000000100000000000010010111111111111111000000000000011010000000000000000000000000001010111111111110101110000000000000010000000000000110011111111110101100000000000010000111111111111100000000000000011111111111111111100000000000001011111111111111011011111111111101001000000000001011111111111111110111111111111111110000000000000011111111111111100001111111111111100111111111111000111111111111111110000000000010000111111111111110100000000000111010000000000000000000000000000001000000000000001001111111111110000111111111111101000000000000010001111111111000110111111111110001100000000000000001111111111111011000000000001011011111111111010001111111111110000000000000001001011111111111100010000000000001000000000000000001000000000000011110000000000010001000000000001110011111111111111001111111111111011000000000000011111111111111111100000000000110011000000000000111100000000000101100000000000111101111111111111100111111111111100100000000000001011000000000000001000000000000000001111111111110010111111111111111011111111111001001111111111111110111111111111111011111111111110100000000000001101000000000000001011111111111111111111111111111010000000000001000000000000000000010000000000001111000000000001010011111111111111100000000000000000000000000000000000000000000101011111111111111001111111111111111000000000000011001111111111110101000000000000000000000000000010001111111111001110000000000001010000000000000000001111111111101001000000000000011111111111110100000000000000000100000000000000010000000000000100100000000000101000000000000001000000000000000011010000000000001001000000000001000000000000000100001111111111101010000000000001000000000000000110101111111111110010000000000000100100000000000101011111111111111110111111111110100100000000000110011111111111111000000000000000101100000000000010011111111111101111000000000000001000000000000000101111111111101111111111111111110011111111111110101111111111111100000000000000100011111111111111010000000000000001000000000000000111111111111101110000000000000001111111111111011100000000000001100000000000000010111111111111111011111111111011100000000000001010000000000000111100000000000011001111111111011100111111111111111011111111111010100000000000000001111111111111100011111111110111011111111111010111111111111111000111111111110111110000000000001100111111111100111111111111111101110000000000000000000000000000001011111111111010011111111111101000111111111111010111111111111101011111111111111001111111111110110111111111111001100000000000000100111111111111111100000000000101100000000000000001000000000000110111111111111110010000000000001100111111111111111011111111111101110000000000000111000000000000001000000000000000000000000000000011000000000000111011111111111101100000000000000101000000000000101100000000000001111111111111111011111111111110011011111111111110000000000000010000111111111101110100000000000001001111111111111100000000000001000100000000000001011111111111101010000000000000100100000000000011000000000000001000000000000010010100000000000000011111111111100101000000000010000011111111111111011111111111101100000000000000001011111111111111010000000000001111000000000001010111111111111101111111111111110010000000000000000111111111111110000000000000001101111111111111100000000000000010100000000000011000000000000000001100000000000101111111111111110101000000000000000100000000000010111111111111111001000000000000111000000000000100000000000000000001000000000000100100000000000001010000000000011000111111111110110011111111111100001111111111101011000000000001001100000000000010010000000000100110000000000001000000000000000010010000000000001101111111111111100111111111111010101111111111001111000000000000010000000000000010010000000000011111000000000010010100000000000111000000000000100010111111111110001011111111111000101111111111010100000000000000101100000000000001101111111111110101000000000001001100000000000000001111111111111101111111111111110111111111111100111111111111101101111111111110001100000000000001100000000000010001000000000000101111111111111110111111111111011101000000000000011111111111111010011111111111101100000000000000001000000000000100100000000000000000000000000000010111111111111010100000000000000011111111111101101011111111111001101111111111111011111111111111111100000000000011010000000000001111111111111111111100000000000011000000000000010010111111111101011011111111111011101111111111110001000000000000011100000000000111010000000000100000111111111110101011111111111111100000000000001111111111111101110011111111111001111111111111110110000000000000110111111111111101000000000000000101000000000000111100000000000001011111111111110101000000000000110011111111111011000000000000000101000000000000000000000000000010001111111111110101000000000000001000000000000001000000000000000100111111111110111111111111111100011111111111110011000000000000100000000000000000100000000000001010000000000000000011111111111101001111111111110010000000000000101000000000000000001111111111101000000000000000101000000000000001100000000000101001111111111111101100000000000000010000000000000000111111111101110011111111111100001111111111101001111111111111000100000000000001000000000000000001000000000000011000000000000100001111111111111010111111111110101011111111111010001111111111101110000000000000111111111111111111000000000000011111000000000000001011111111111001001111111111111110000000000000000011111111111101111111111111100111000000000001001000000000000000110000000000001000111111111111001011111111111011111111111111111110111111111110001011111111111100111111111111101100000000000001001100000000000001010000000000100000000000000000101100000000000111000000000000010010111111111111100011111111111010111111111111101101111111111111110000000000000101011111111111111011111111111110101011111111111001101111111111101101111111111110011011111111111100001111111111100100000000000000000000000000000011110000000000001010000000000000111111111111111011101111111111110100111111111111111111111111111001000000000000000000111111111111010100000000000001110000000000010110000000000000011011111111111111000000000000001111111111111111011011111111111001101111111111101010111111111110100100000000000111000000000000001001000000000000010100000000000111001111111111111010111111111110010111111111111011011111111111011101000000000001000000000000000110100000000000001110000000000001011000000000000001010000000000001001111111111101111011111111111010111111111111101110111111111111101100000000000100110000000000011101111111111111011111111111111101011111111111111111111111111111110000000000000011011111111111101111000000000000100000000000000000000000000000010101111111111111110100000000000100000000000000000111111111111110010111111111111010101111111111101000111111111111111011111111111111000000000000010110111111111111101011111111111001110000000000000110111111111110101000000000000000111111111111110100000000000000010111111111111011110000000000000110000000000001101100000000000000001111111111101110000000000001011011111111111011111111111111110001111111111111101100000000000110000000000000101010000000000000001011111111111101110000000000001001000000000000111011111111111101101111111111011111000000000000000111111111111100101111111111111001111111111111000011111111111101010000000000011000111111111111100111111111111001100000000000000110000000000000000100000000000011100000000000000101000000000001010111111111111100111111111111010011111111111111100000000000000000000000000000000011000000000000000000000000000000001111111111011010111111111111101000000000000101100000000000000010111111111111100100000000000101010000000000011000000000000001011000000000000011000000000000000111111111111111010000000000000000101111111111111010111111111111011011111111111101100000000000000110000000000000011100000000001001101111111111111110000000000001001011111111111101001111111111111101000000000000001011111111111000101111111111110110111111111101110011111111111101100000000000100001111111111111000111111111111101011111111111110111111111111111100111111111111011011111111111011111111111111111111100000000000000101111111111111101111111111111111100000000000001000000000000000010111111111110111100000000000000000000000000001100000000000000000011111111111000101111111111010100000000000001101011111111111100101111111111001101000000000000111111111111111100000000000000000101000000000000000011111111110111101111111111000001000000000010001100000000000101110000000000000101000000000000101111111111111010000000000000011100000000000000010111111111110111011111111111111010111111111111101100000000000001100000000000001111000000000000101100000000000111010000000000101110000000000001101011111111110111011111111111010100111111111111100111111111111100101111111111101111000000000000111000000000000000100000000000100000111111111110110111111111111010001111111111100111000000000000010100000000000010010000000000011011000000000000001000000000000011010000000000010010000000000010101000000000000001011111111111100010111111111111110011111111111010000000000000010010000000000000010000000000000011000000000000101010000000000000101111111111111100000000000000000111111111111110101011111111111101100000000000010010111111111110101111111111111101001111111111110110111111111101111111111111110101111111111110100110000000000010100100000000000001111111111111010101111111111111111100000000000101000000000000110100000000000001111100000000000000011111111111110010000000000010101111111111111101101111111111110000000000000001101011111111111010000000000000000110111111111111001100000000000110010000000000000101111111111111100011111111111101010000000000001111000000000000011111111111111100011111111111100011000000000001001000000000000000000000000000000101000000000000010111111111111111101111111111101011000000000000000011111111111010100000000000001110111111111111100011111111111100101111111111111110000000000000001000000000000000101111111111100111000000000000101100000000000011000000000000001100111111111110110111111111111001000000000000000110000000000001011000000000000111010000000000010100000000000000111100000000000110000000000000010100111111111111010111111111111001010000000000100011000000000000001011111111111010111111111111110010000000000000011000000000000110011111111111100011111111111111111100000000000010010000000000011111000000000000100011111111111111110000000000000000000000000000101111111111111000001111111111011101000000000001001111111111110110001111111111111111000000000000010100000000000101010000000000010101111111111111010111111111111001100000000000010100111111111111100000000000000010101111111111110101000000000001100111111111111011011111111111101000111111111111101000000000000101100000000000100111000000000001100100000000000100010000000000001110111111111110100100000000000000101111111111111011111111111111110000000000000000001111111111111000111111111110100011111111111001100000000000000100000000000001010100000000000000001111111111111101000000000001011000000000000100000000000000000000111111111111111111111111111110001111111111110011111111111110000100000000000110110000000000011110000000000000000011111111111010000000000000000010000000000001101100000000000001010000000000010111111111111111110111111111111001000000000000001000111111111110101000000000000010001111111111111111000000000001010011111111111110100000000000100010000000000000000011111111111110001111111111111100111111111101100011111111111100111111111111101111000000000000011011111111111100011111111111011000111111111110111011111111111010101111111111111010111111111110011000000000000000000000000000110100000000000000000000000000000010001111111111111001111111111111010000000000000001010000000000000110000000000000100100000000000011101111111111111110000000000000011111111111111101111111111111111011111111111111101000000000000000000000000000000000000000000001000100000000001000000000000000001000000000000000001111111111111010101111111111010111111111111111001100000000001000100000000000100001111111111110011011111111111111001111111111110111000000000000100011111111111000111111111111011111000000000000001111111111111111011111111111101010111111111111100111111111111001001111111111100110000000000000011111111111111100001111111111110001000000000001001000000000000101011111111111101011111111111110101111111111110110011111111111101100111111111111010111111111111110100000000000000000000000000001000100000000000101000000000000001100000000000001000000000000000011111111111111100110111111111111000000000000000101010000000000111010111111111111011100000000000010000000000000010011111111111111001100000000000101110000000000001011111111111111100111111111111110000000000000001000111111111111101011111111111011101111111111111110111111111110110011111111111110111111111111111011111111111111010111111111110011111111111111101100000000000010000000000000001101000000000000110011111111111110011011111111111111000000000000001110111111111111100111111111111100010000000000010010111111111101011111111111111000000000000000010101111111111110101100000000000010000000000000000011000000000000110011111111111110100000000000000010000000000000000111111111110111011111111111100001000000000000110111111111111011100000000000001001111111111111001111111111111101010000000000100011000000000001001000000000000000111111111111111101111111111111011011111111111111111111111111111101000000000000010100000000000011110000000000100101000000000001010111111111111111001111111111110001111111111111011011111111111100011111111111110101000000000000000011111111111111001111111111010011111111111110100111111111111101101111111111100111000000000000011111111111111101110000000000001111000000000001001011111111110010001111111111010111000000000010010100000000000000011111111111111100000000000010011100000000000100110000000000011000000000000010011100000000000100101111111111111100000000000000101011111111111110011111111111100001111111111111111100000000000000000000000000001000000000000001010000000000000011010000000000000001000000000000110100000000001101100000000000001011000000000000000111111111111011111111111111100100000000000001000100000000000110110000000000010100111111111111100000000000000101011111111111001101000000000000101011111111110111101111111111101110000000000001000111111111111110101111111111111010000000000001001111111111111111011111111111110111000000000011001100000000001101010000000000011101000000000000000111111111111110011111111111110000000000000001000100000000000000111111111111100110000000000000000011111111111101111111111111111000111111111111111000000000000010111111111111110001111111111101100011111111111011100000000000001100111111111110110111111111110110111111111111011111000000000000100111111111111110011111111111111010111111111111010111111111111010111111111111111100111111111111111011111111111000101111111111110011000000000000111011111111111110100000000000000101000000000000010100000000000100100000000000001111111111111111100100000000000001001111111111101010000000000001011100000000000111000000000000000010000000000000101000000000000100000000000000100101000000000001100000000000000000000000000000011001111111111111101100000000000001111111111111110010111111111111101000000000000000010000000000010101000000000000001011111111111011100000000000000101111111111111110011111111111101001111111111101100000000000000111011111111111100010000000000000111000000000001001111111111111110100000000000001111111111111111111100000000000000111111111111101100111111111111010011111111111100000000000000001010000000000000000011111111110100111111111111100100000000000010000000000000000111001111111111101001000000000000000111111111111001100000000000001000000000000001010000000000000101010000000000001111000000000000111011111111111011011111111111111110000000000000000011111111111011000000000000001110000000000010101011111111111111101111111111111110111111111110110000000000000101001111111111110110111111111110011111111111111111111111111111110010111111111110100111111111111101001111111111100000111111111111111011111111111110101111111111111100000000000000000100000000000110110000000000011110111111111110111011111111111100001111111111001110000000000001000100000000000001101111111111101100000000000000110100000000000000001111111111110111000000000010001000000000001010100000000000010101111111111111011111111111111110001111111111100000111111111111011011111111111001010000000000000010111111111100010011111111111001101111111111011110111111111111101000000000000011001111111111110101000000000000000111111111111100110000000000011010111111111111011011111111111100011111111111011111111111111111011111111111111110110000000000001010000000000001011111111111111100101111111111100111000000000000101000000000000001000000000000000000000000000001010100000000000100101111111111110010111111111111100000000000000001100000000000000000000000000000101111111111111101101111111111110001000000000010011000000000000011000000000000100101000000000000001100000000000000010000000000011110111111111101111011111111111011111111111111011000000000000001000000000000000110001111111111110110000000000010001111111111111111000000000000000000000000000000011011111111111110101111111111111000000000000001101100000000000110101111111111100111000000000001111111111111111100101111111111001101000000000000100100000000000000101111111111110101000000000000000011111111111100000000000000000011000000000000011000000000000000000000000000010001000000000000100000000000000100001111111111110001111111111110110100000000000001010000000000000101000000000000000011111111111111001111111111101011111111111111100000000000000011010000000000000100111111111101110000000000000010010000000000000001000000000010010000000000000000110000000000000000111111111110000000000000000011000000000000001001111111111111000011111111111001110000000000001000000000000001000011111111111110111111111111110100000000000000100111111111111111111111111111111100000000000000000100000000000100000000000000000000111111111110111111111111111100011111111111111010111111111111101000000000000001000000000000000000000000000000000000000000000001001111111111110100111111111110110011111111111101000000000000010001111111111111000000000000000010001111111111111101111111111111011000000000000001011111111111111101111111111111111011111111111011111111111111100110000000000000000111111111111100101111111111110110111111111111011111111111111111110000000000001100000000000000000100000000000000101111111111110111000000000000110111111111111111000000000000000011000000000001010000000000000000100000000000010010000000000000010000000000000001111111111111101110111111111111111111111111110111101111111111111011111111111111101100000000000011001111111111111100000000000000111111111111111110011111111111111101000000000000000000000000000000101111111111111000000000000001111000000000000100010000000000000100000000000000000000000000000000000000000000000000000000000000010000000000000010000000000000000011111111111111101000000000000000100000000000000110111111111111101011111111111101000000000000001011111111111111011100000000000000010000000000001111111111111111000111111111111111111111111111111101111111111111000111111111111110010000000000000011111111111111101011111111111101001111111111110111000000000000000111111111111101011111111111111001111111111111100100000000000001100000000000000100000000000000011111111111111101101111111111110111000000000000000000000000000000010000000000010011111111111111011000000000000000100000000000000010000000000000111100000000000000111111111111111111111111111111110100000000000001001111111111101110111111111111000100000000000010000000000000001010000000000000100011111111111111110000000000000000000000000000010100000000000001001111111111111010000000000000101011111111111110010000000000010100000000000000000111111111111111101111111111111101000000000000010011111111111101111111111111111010111111111111001111111111111101000000000000000001111111111111011011111111111111111111111111101101111111111111100000000000000100110000000000001011111111111111111111111111111010101111111111111010111111111111110011111111111110110000000000001000111111111111111111111111111101001111111111111111000000000000101011111111111010000000000000000010000000000000001100000000000010010000000000010010000000000000111111111111111110111111111111111110111111111111011000000000000011001111111111111011000000000001011000000000000010111111111111111111111111111111101011111111111110111111111111100101000000000000010000000000000001110000000000011101000000000000011000000000000000011111111111110010000000000001001100000000000011000000000000001000111111111111101011111111111101001111111111111101111111111111000011111111111101100000000000000000111111111111100100000000000000001111111111100000000000000000001000000000000001101111111111101011000000000000000011111111111110110000000000000110111111111110101100000000000011101111111111111111000000000000011100000000000001010000000000000000000000000001001100000000000000110000000000010001111111111110000011111111110010111111111110110010000000000000111111111111111011100000000001000101111111111111110111111111111010000000000000101010000000000001011000000000000000110000000000000101111111111101111111111111111001100000000000110000111111111110011100000000000101010000000000100000000000000001001000000000000010011111111111101010111111111111000011111111111010101111111111110110111111111110101011111111111110011111111111011010111111111101110011111111111001011111111111110001111111111110101100000000001100000000000000000100000000000000100000000000000010110000000000001110000000000001111000000000000011111111111111100011000000000000011011111111111111101111111111011101000000000001010111111111111111010000000000010111000000000011001111111111111011101111111111110011000000000000101011111111111100000000000000011101111111111110101011111111111100000000000000100000111111111110100111111111110100001111111111110101111111111110110000000000000011000000000000101100111111111111011111111111111111110000000000011011000000000011100100000000000001011111111111011101000000000000000111111111110010101111111111110011111111111111101011111111111001011111111111110101000000000001001100000000000000100000000000000001111111111111100000000000000000101111111111111100111111111111101011111111111111110000000000000000000000000000010000000000000100001111111111101011000000000010000000000000000011101111111111000110000000000000101011111111110111011111111111010100000000000000100000000000000010110000000000010100000000000000101000000000000010000000000000000000111111111111111011111111111111100000000000011011000000000010011011111111111101101111111111000001000000000001010000000000000000001111111111000011000000000001001100000000001011101111111111100000000000000001001000000000000010001111111111001111000000000010011011111111111101101111111110110101000000000000101011111111111001011111111111100000000000000000011011111111110110011111111111100101111111111111110011111111111010111111111111100100000000000010001000000000000000110000000000011101000000000001110011111111111111001111111111111000111111111111110111111111111110100000000000000110111111111111000000000000000100010000000000000011000000000000110100000000000000101111111111110101111111111110111011111111111010101111111111011101111111111111100100000000000010111111111111111100000000000000100111111111111110001111111111111010000000000010001100000000001011000000000000000000000000000010010000000000001000001111111111100100000000000001110111111111111000111111111111011011000000000000111111111111111110011111111111100110111111111111010111111111111110111111111111110111000000000001000000000000001011001111111111110010111111111110010111111111111111000000000000010111111111111111010000000000000100001111111111111010000000000000100011111111111111001111111111111011000000000000001000000000000000111111111111110001111111111110010011111111111011001111111111111000000000000000100000000000000111110000000000110101000000000001000111111111111010101111111111101111000000000010111011111111111000110000000000001100000000000000010011111111110111101111111111101111000000000000011111111111111000010000000000001011000000000000010111111111110100100000000000011100000000000001110011111111111111101111111111011110111111111110010111111111111101010000000000100101000000000000101000000000000101000000000000001111000000000000000000000000000011001111111111110100111111111111111100000000000010111111111111101110111111111111101100000000000100100000000000000110111111111111110111111111111011010000000000001100000000000000111100000000000001000000000000000101111111111111101000000000000001000000000000001010000000000000100011111111111111011111111111100001000000000010111000000000000001011111111111011001000000000000111111111111111101111111111111101011111111111111000111111111111011001111111111101010111111111111010111111111111101001111111111111000000000000000000000000000000001000000000000010011111111111111110111111111111001111111111111101010000000000001010011111111111100110000000000000011111111111111110100000000000010001111111111110011111111111110111011111111111111110000000000010010111111111110111011111111111101100000000000001011111111111110100011111111111111111111111111110001111111111111110111111111111101011111111111111110111111111111001011111111111111011111111111111011000000000000001100000000000010111111111111111100111111111111111000000000000011101111111111110101000000000000101000000000000000100000000000000110000000000000001000000000000001100000000000011000111111111111001000000000000000001111111111111111111111111101110100000000000000000000000000011011111111111111110100000000000110001111111111011110111111111110010000000000000001111111111111100110111111111111101000000000000001000000000000000011000000000000100011111111111101100000000000011100111111111110111111111111111100111111111111110100000000000000001011111111111011101111111111110101111111111111100000000000000100111111111111110111111111111111000100000000000111001111111111111011000000000000001111111111111111100000000000000001111111111111000011111111111001011111111111110010000000000000010100000000001111010000000000111110111111111111011100000000000011010000000000001110000000000001000000000000000100100000000000000010000000000000000011111111111101110000000000100101111111111111000100000000000010101111111111110011111111111111100111111111111111111111111111111101111111111110011100000000000011100000000000011010111111111110111100000000000000000000000000000000111111111111100011111111111111000000000000001011111111111101101011111111110100101111111111100001111111111111010111111111111000001111111111111110111111111110010111111111111010100000000000010010000000000000011000000000000000000000000000000000111111111110001011111111111101111111111111101001111111111110000111111111111011011111111111101111111111111111111100000000000010111111111111110100000000000000001111111111111010101111111111100011111111111111010000000000000001011111111111101011111111111110000111111111110111011111111111101000111111111111011011111111111010111111111111110010000000000000001011111111111100001111111111101111000000000001001000000000000001100000000000011000000000000001000100000000000000111111111111101111111111111111101100000000000001100000000000001001111111111111001000000000000010000000000000000010111111111111000111111111111101010000000000001001111111111111010011111111111110110000000000010010000000000000011111111111111111011111111111101010111111111111010000000000000101100000000000000001111111111111011100000000001001000000000000001101111111111111101000000000000111010000000000011001111111111111100011111111111111100000000000001111000000000001011011111111111100100000000000000001000000000000101111111111111110001111111111110011000000000001011100000000000011101111111111110001000000000000001000000000000001101111111111010111000000000000011100000000000010100000000000001111000000000000100000000000000100001111111111111111000000000001110100000000000100110000000000000000000000000001110011111111111011011111111111110011000000000010000000000000000000011111111111110011111111111111101111111111111011001111111111101001111111111110110111111111111011111111111111001010111111111111011011111111111111011111111111010101000000000001100111111111111111011111111111101100000000000001010000000000000000000000000000001100000000000000111100000000001001110000000000001101000000000000010100000000000110110000000000011111000000000000011000000000000001111111111111111001111111111111111000000000000010100000000000000111000000000000000011111111111010100000000000001001111111111110101111111111111011001111111111110010111111111101110100000000000010101111111111101101000000000010010100000000000000111111111111111001000000000001001000000000000010001111111111110101000000000000111111111111111111000000000000011110000000000000011100000000000011000000000000000101000000000001100100000000000010000000000000000000000000000001000100000000000101110000000000000111000000000000000000000000000001100000000000010100000000000001000011111111111101100000000000000010000000000001101100000000000110110000000000000101111111111111101100000000000001100000000000000011111111111111111111111111111101001111111111101100111111111111101011111111111110011111111111101111111111111111001111111111111110001111111111110000111111111110110100000000001011010000000000110011111111111110110000000000000010100000000000001111000000000001000000000000000111010000000000001100111111111110101111111111111000001111111111111100000000000000010100000000000100111111111111100100000000000001010011111111111101100000000000000001111111111111001011111111111100110000000000010101000000000000010100000000000001000000000000000011000000000010111100000000000111011111111111110000111111111111000000000000001000100000000000001110111111111111011000000000001000000000000000001101000000000000010000000000000111000000000000001001111111111111011111111111111010101111111111111010111111111111010100000000000000001111111111110101000000000001110100000000000001001111111111111110000000000001010011111111111101100000000000000011111111111111010111111111111111001111111111111100000000000000000100000000000110010000000000000010000000000000010100000000000001001111111111011101111111111111000100000000000010010000000000000001111111111111110111111111111110100000000000001001000000000000000011111111111011001111111111010001111111111111111111111111111010111111111111101110111111111111111011111111111110010000000000010011000000000000111100000000000001000000000000001011000000000000110111111111111100000000000000000000111111111111110111111111111101010000000000001010111111111111001111111111111111101111111111100110000000000000010000000000000001001111111111110101000000000000000011111111111011011111111111110111000000000000000100000000000001100000000000000110000000000000010111111111111111110000000000001110111111111111010100000000000011000000000000001010000000000000110011111111111011101111111111100110111111111111111111111111110111101111111111100011000000000001011011111111111111110000000000011100000000000000000111111111111111010000000000001100111111111111110000000000000000110000000000000111000000000000011111111111111111111111111111010000111111111110011111111111111100111111111110110100000000000000111111111111111011101111111111000100000000000000000000000000000011001111111111001001000000000000000000000000000011100000000000001101000000000010111100000000000010111111111111110010111111111111000111111111111010101111111111110010111111111111001011111111111101000000000000011101111111111100011111111111111101100000000000100001111111111111000100000000000100010000000000011111111111111111010111111111111101001111111111110000000000000000100011111111111001000000000000101101111111111101100111111111111011100000000000001101111111111111100000000000000011011111111111111111111111111111101000000000000101000000000000010100111111111111111000000000000111010000000000010111111111111111001111111111111100000000000000001100111111111111001100000000000111100000000000011010111111111110111100000000000110000000000000011110000000000000010100000000000100011111111111011101000000000000001111111111110111111111111111111001111111111110100011111111110111100000000000001011111111111111101011111111111111000000000000010101111111111111011100000000000010110000000000000110111111111111100100000000000100010000000000001011000000000000110011111111111011110000000000110001111111111111001000000000000101100000000000111010000000000000000100000000001000110000000000011100111111111110110100000000000100011111111111110001111111111111111111111111111011001111111111111001000000000001010111111111111111111111111111100101111111111111111011111111111101010000000000001100000000000000001000000000000010111111111111111100000000000001010011111111111111000000000000000100000000000000010100000000000001100000000000100000111111111110101000000000000001001111111111101111111111111111001000000000000000100000000000001000111111111111101011111111111000001111111111101011111111111111101011111111110111111111111111101101111111111110110011111111111001110000000000000101000000000000100100000000010000110000000000011101000000000000001000000000000001101111111111101001111111111111111100000000000001110000000000000000111111111111100100000000000111110000000000010011000000000000101100000000000001000000000000001011111111111111100000000000000000000000000000001101000000000000000000000000000011011111111111110001111111111110001111111111111011011111111111110001111111111111101111111111110100101111111111111010111111111110111000000000000010010000000000000010111111111110011011111111111111101111111111101101000000000000010000000000000001011111111111101011111111111111011100000000000000011111111111111010111111111111000011111111110110100000000000001110000000000000000111111111111101011111111111110001111111111100100011111111111011100000000000000100111111111101101100000000000010101111111111111100111111111110001000000000000000000000000000010010111111111110010100000000000100100000000000100010111111111110010100000000000000111111111111111001111111111111110011111111111101001111111111101110111111111111011011111111111111010000000000000110111111111111001011111111111101100000000000111110111111111110110000000000000001110000000000011100111111111101101000000000000010100000000000010111111111111111000100000000000000001111111111110110111111111111010100000000000011010000000000000100111111111110100100000000000000010000000000000000000000000000101111111111111100111111111111101101000000000001000011111111111100000000000000000010000000000000001100000000000011011111111111110110000000000000100000000000000000101111111111011100000000000000010011111111111100001111111111111111000000000000010011111111111010100000000000000110111111111101110011111111111000110000000000100100111111111110101111111111110110010000000000010011000000000000000000000000000110001111111111110100111111111111110100000000000100010000000000000111111111111111011111111111111110011111111111111111111111111110100011111111111111011111111111100111111111111110101100000000000000100000000000001001000000000001011000000000000001001111111111110111000000000000010100000000000100000000000000011100000000000001010011111111111100100000000000000111111111111110011111111111111110011111111111110111111111111111110000000000000111101111111111110101000000000000010100000000000011010000000000000001000000000000010000000000000001100000000000011001000000000000011100000000000010001111111111101100111111111110101011111111110111111111111111101011111111111111110100000000000000111111111111110001111111111111011111111111111010001111111111101101000000000000000011111111111011100000000000000101000000000010010000000000000011000000000000001010111111111110111011111111111011001111111111111100000000000000011011111111111100000000000000010000000000000000011111111111111101110000000000001101111111111111011111111111111101011111111111010111111111111111000111111111111111001111111111110011111111111111111100000000001010101111111111101111000000000001101100000000001000000000000000011110111111111111110100000000000011000000000000001001111111111111100100000000000010000000000000001110000000000000001100000000000000000000000000010011111111111111100011111111111101010000000000000101111111111111101100000000000100100000000000000101111111111111110111111111111110110000000000000111111111111110111100000000000000100000000000001011000000000010001000000000000111100000000000011100111111111110001011111111111100011111111111101001111111111111011011111111111011101111111111111000000000000000110100000000000001110000000000000110000000000000010011111111111100001111111111100111111111111111010011111111111110110000000000000011000000000000101100000000000110000000000000011101000000000000010000000000000000000000000000000001111111111111111111111111111101111111111111111001111111111111110000000000000011010000000000110001111111111111110111111111111111011111111111101111111111111110100111111111111110110000000000001110111111111111110100000000000000110000000000000000111111111111100111111111111101000000000000010011000000000000001011111111111101100000000000001000000000000000011011111111111111001111111111110101000000000001001100000000000010110000000000001111000000000000110000000000000010000000000000011111111111111111001100000000000000100000000000000011000000000001110100000000001001000000000000000100111111111111110111111111111010011111111111100111111111111111101000000000000000110000000000000001111111111110101100000000000010000000000000000010111111111111111111111111111011001111111111111011111111111111011100000000000001010000000000000111111111111110110111111111111011011111111111110010111111111110111111111111111011101111111111011001000000000000010000000000000000111111111111110101111111111110101100000000000000000000000000000100000000000000010000000000000011001111111111101110000000000000000000000000000000100000000000000110000000000000000000000000000101100000000000000010000000000001100000000000000110010000000000010110111111111111001100000000000001010000000000000100111111111111001011111111111111100000000000010000111111111111101011111111111011011111111111100011000000000000100000000000000110010000000000010100000000000000100000000000000000111111111111110010111111111111101111111111111010001111111111110001000000000000011111111111111000101111111111111000000000000000100000000000000001101111111111100011000000000000000111111111111110000000000000000110111111111111110000000000000011000000000000010010000000000000000111111111111011111111111111111110000000000000001011111111111000111111111111001100000000000000111011111111111110100000000000001110111111111111101011111111110100001111111110101001111111111111111111111111111110011111111111111011000000000000100000000000000010100000000000010100111111111111111000000000000000010000000000000111111111111110110100000000000011101111111111111000000000000000000111111111111100101111111111101110000000000000101000000000000001110000000000001001111111111111010100000000000010000000000000001110000000000001000000000000000010100000000000001100000000000001011100000000000000000000000000000001000000000000100000000000000011110000000000010010000000000001001000000000000101000000000000000101111111111111010011111111110110011111111111011011111111111111000011111111111111010000000000011110000000000010000100000000001001110000000000001101000000000000000011111111111000001111111111011101000000000000011000000000000010100000000000001001000000000010110100000000000011100000000000001101111111111111010011111111111011111111111111010001111111111100110111111111110011001111111111100100111111111110011000000000000000000000000000001101000000000000000011111111111100011111111111111010000000000000011011111111111111111111111111110100000000000000110000000000000001100000000000000000000000000010001000000000000010110000000000001001000000000000010000000000000001011111111111111110111111111111011000000000000011100000000000011110111111111111110011111111111110110000000000011110000000000000111000000000000010000000000000010110000000000010010100000000000001111111111111111011000000000001011111111111111111001111111111110111000000000000100000000000000000101111111111101011000000000000100111111111111011101111111111111010000000000001011011111111111110101111111111011111111111111111000100000000000010100000000000000100111111111111110100000000000001001111111111101000000000000010101100000000000111010000000000100000000000000001100000000000000100000000000000000000000000000000100011111111111111011111111111110000111111111101000011111111111000011111111111110001000000000000110000000000000001110000000000000001000000000010011100000000000011110000000000000000111111111111110100000000000001010000000000001100000000000000011000000000000110100000000000001011111111111110111111111111111011111111111111110101111111111111111011111111111110000000000000010110111111111101011000000000000011010000000000101011000000000000100000000000000000101111111111101011000000000000010100000000000010010000000000000101111111111110011111111111111100001111111111111111000000000001001100000000000000010000000000010111000000000001110100000000000000000000000000001010000000000001111000000000000010000000000000010100000000000001100000000000000011101111111111111110111111111111101011111111110110011111111111010111000000000000101100000000000000001111111111111111000000000000101000000000000101101111111111101100111111111111101011111111111101011111111111011000000000000000010100000000000100100000000000001110111111111111110111111111111100101111111111011111000000000010110100000000000101001111111111100111000000000001000111111111111101011111111111100100000000000001110011111111111110000000000000010011000000000000100011111111111100101111111111110011000000000001010000000000000011001111111111111110111111111111101100000000000010100000000000000111111111111111101011111111111010111111111111110101000000000000011011111111111011111111111111111100000000000001100000000000000000000000000000010000111111111100000011111111111010011111111111110111111111111111110111111111111110010000000000010000000000000001110100000000000111110000000000011000111111111110011011111111110111111111111111101001000000000000010100000000000001000000000000100110000000000010011100000000000101000000000000010110000000000000010011111111111101101111111111111011000000000000000111111111110100001111111111100001000000000000011011111111111110111111111111110100000000000000001000000000000010000000000000001001000000000000000100000000000000011111111111101110000000000000110111111111111110110000000000000010111111111111101100000000000111100000000000100010000000000001000000000000000000110000000000000000111111111111100011111111111011101111111111010101111111111110111011111111111111001111111111111100000000000001001100000000000001001111111111110110000000000010001100000000000000011111111111110100111111111100011011111111110110011111111111111000000000000001000011111111111111010000000000000100000000000001110000000000000111000000000000000100111111111110011111111111111011111111111111110000000000000001010011111111111011110000000000010101000000000001101100000000000111110000000000011001000000000000011111111111111010110000000000000010000000000001011011111111111101011111111111111001111111111111011111111111111101000000000000000000000000000001000100000000000000001111111111100011000000000000000111111111111100111111111111001001000000000000010111111111111100110000000000000000111111111110011100000000000011110000000000011101111111111111101000000000000000111111111111111010111111111111100011111111111000100000000000000011000000000001100100000000000110000000000000000010111111111111110000000000000001011111111111111011000000000001010100000000000010001111111111111101111111111111010100000000000001001111111111110000111111111111010111111111111100101111111111110001000000000000011000000000000001111111111111110001000000000000101000000000000101110000000000000110111111111111011000000000000001000000000000001101111111111110100000000000000010101111111111111111111111111110001011111111111100001111111111111001000000000000101000000000000000011111111111111000000000000000010000000000000100001111111111100001000000000001100011111111111111011111111111111101111111111111111111111111111100011111111111110100111111111111000111111111111110111111111111100010000000000001011000000000000001110000000000010100111111111111111000000000000010011111111111111111111111111101111111111111111000000000000000010010111111111100000111111111111011011111111111001100111111111111110111111111111000001111111111100010000000000000011011111111111011111111111111001100111111111110100100000000000100010000000000010001111111111111110011111111111110110000000000010001000000000000001100000000000011010000000000001010111111111111011111111111111111101111111111101001000000000000101011111111111110001111111111111001000000000001111100000000000011010000000000000110000000000001011011111111111000010000000000000010000000000000100100000000000101000000000000010001111111111100110111111111111101000000000000010000000000000001110000000000000110101111111111110110111111111110101000000000000010110000000000000111000000000000001000000000000101010000000000010100000000000000010100000000000100111111111111110111111111111110000111111111111110000000000000000110000000000001000000000000000110010000000000010111111111111111011011111111111010111111111111110111000000000000101011111111111101000000000000000000000000000000101100000000000110011111111111111010000000000001110000000000000011110000000000001111111111111111001111111111111110011111111111101001111111111110110111111111111000011111111111100101000000000001001000000000000110000000000000001111000000000000000011111111111101111111111111110101000000000000000000000000001000000000000000001100111111111111001000000000000000110000000000101001111111111110010011111111111011010000000000000101111111111101001011111111111000001111111111100111000000000001010011111111111011111111111111100111000000000001010111111111111111000000000000000000000000000000010000000000000001001111111111101100000000000010011000000000000000000000000000011100111111111110111100000000000000111111111111111001111111111111110100000000000100010000000000100100000000000001101011111111111111110000000000011010111111111110110011111111111110011111111111110111111111111101111011111111110110110000000000000101000000000000101000000000001000011111111111111001111111111110110011111111111000011111111111011110111111111110111111111111111001100000000000001000111111111111101100000000001000100000000000110000000000000000100100000000000101000000000000011011111111111011100111111111110000101111111111001100000000000000111000000000000000110000000000010010111111111111101011111111111110011111111111111101000000000001000100000000000110011111111111110011111111111111110011111111110100101111111111010100111111111110000111111111111110001111111111110111111111111110101011111111111010001111111111110000000000000001110000000000000000000000000000100000111111111111000111111111111101010000000000001010000000000000001100000000000011000000000000010101111111111111101111111111111000010000000000010101000000000000110111111111111100001111111111010101000000000001110100000000000001101111111111011101111111111111101011111111111100011111111111110001000000000000000011111111111001011111111111100111000000000000111100000000000001110000000000001010000000000000110111111111111110001111111111111111000000000000010000000000000010000000000000001111000000000000100100000000000010110000000000001001000000000001100100000000000010110000000000001001111111111110100011111111110111001111111111111010111111111110001000000000000000000000000000100100111111111111000100000000000000101111111111111001111111111110011111111111111000100000000000001010111111111110111111111111111000011111111111101111000000000001100000000000000001001111111111110111000000000010010100000000000010100000000000001100000000000001001100000000000110000000000000001111000000000001111011111111111110001111111111010011111111111110001111111111111101011111111111110000111111111101010111111111111000011111111111111101000000000000101111111111111111001111111111110011111111111110000111111111111010011111111111101010000000000000100111111111111101101111111111110111000000000001010111111111111101011111111111101101111111111111001111111111111001011111111111111110111111111110011011111111111010111111111111111010111111111111111100000000000011110000000000001001000000000000011100000000000001110000000000000011000000000010001000000000001010010000000000000101111111111110101000000000000000110000000000000111000000000000000011111111111010000000000000010010000000000000110111111111110111100000000000000001000000000001101011111111111111011111111111110111111111111111101000000000000010111111111111111010000000000000011111111111111111011111111111100100000000000001110000000000000011011111111111101000000000000000010000000000000001111111111111110000000000000000000011111111111100001111111111110110111111111110111111111111111100011111111111101110000000000000100111111111111101001111111111101101000000000000010000000000000001101111111111100100000000000000100100000000000011000000000000000001111111111111001111111111111010101111111111110101111111111110111011111111111010100000000000001010000000000000110000000000000100000000000000010101000000000010000100000000000010111111111111111011000000000000110000000000000001100000000000001001000000000000111000000000000011100000000000000000000000000000011111111111111011011111111111110000000000000001011000000000000010111111111111101111111111111111010011111111111000101111111111011000111111111111100100000000000011110000000000010101111111111110111011111111111111100000000000011001000000000000000011111111111110000000000000001011111111111111110100000000000000000000000000001110000000000000110100000000000010100000000000001111000000000000011011111111110111111111111111110001000000000000001011111111111111001111111111110000111111111111111100000000000011001111111111110100000000000000000011111111111000100000000000000011111111111110110000000000000000011111111111100111111111111111111011111111111110011111111111101100000000000000100111111111111110100000000000000100000000000001000100000000000010111111111111110010000000000000101011111111111011100000000000001001000000000001100000000000000000011111111111101010000000000010110100000000000111110000000000001101000000000001011000000000000001010000000000010100111111111111100111111111110111011111111111001000000000000001011100000000000010110000000000000001111111111110100100000000000000100000000000001010111111111111000011111111110110111111111111101011111111111110110000000000000000101111111111111000000000000000000000000000000001000000000000101010000000000001100011111111111110101111111111111001000000000000010100000000000010000000000000001010000000000001010000000000000100010000000000011101111111111110111111111111110111111111111111100000111111111111101000000000000011000000000000000100000000000001000000000000000010100000000000010111000000000001100100000000000100001111111111110001000000000000100000000000000100111111111111111011111111111111100111111111111100001111111111110111111111111111100100000000000011010000000000000100000000000000100111111111111110010000000000000000000000000001001100000000000000110000000000010001111111111110111011111111110100111111111111011010000000000010111100000000000000101111111111111110000000000000000000000000000101100000000000000111000000000001101111111111111010011111111111101111000000000001100000000000000111110000000000001110000000000000111100000000000101000000000000001000111111111111110111111111111011011111111111111010111111111110110111111111111001110000000000000001000000000000101111111111111100011111111111101110111111111111011011111111111101000000000000000011000000000001010100000000000011100000000000011111000000000000000000000000000110110000000000001001111111111111000111111111111111111111111111110110111111111111110111111111111100111111111111101110000000000001111100000000000100000000000000000110111111111100100011111111110000001111111111011000111111111110101000000000000000011111111111011011000000000000011111111111111111100000000000010000111111111101111011111111110111111111111111110000000000000000000111111111111010101111111111100010000000000011001100000000000100111111111111011001111111111101111011111111111100011111111111110100111111111111110011111111111010011111111111111011000000000000101011111111111011001111111111110110111111111111100011111111111010100000000000000111000000000001010011111111111011001111111111101001000000000000000011111111111000001111111111111011000000000001111111111111111111101111111111001011000000000001101111111111111001011111111111100111000000000000111011111111111011001111111111010011111111111110100000000000000000000000000000000000111111111110011000000000000011100000000000010011111111111111010111111111111101010000000000001001000000000000101111111111111100101111111111111101111111111111101111111111111010001111111111111100111111111111110111111111111011010000000000011100000000000000110000000000000011100000000000010000000000000000101000000000000100000000000000000110111111111111100111111111111110111111111111111000111111111110001000000000000000110000000000000001111111111110110011111111111101111111111111110100111111111101101011111111111110010000000000000110000000000000000011111111111110001111111111111001000000000000000011111111111101111111111111100100111111111111000111111111111101000000000000001100111111111111100000000000000010000000000000001001000000000000111000000000000100100000000000000000000000000000101100000000000011110000000000001010111111111111101000000000000000000000000000000000111111111111111111111111111111001111111111110100000000000000001011111111111101110000000000000101111111111110011111111111110011111111111111111111000000000000101011111111111011110000000000001001000000000000010111111111111100000000000000011011111111111111100000000000000100111111111111111111111111111111110000000000000010011111111111110001111111111111110011111111111010001111111111110111000000000101011000000000001001100000000000010101000000000011011000000000001001001111111111111110000000000000011100000000000001111111111111110010000000000000000000000000000010110000000000011111000000000001011100000000000111010000000000010101000000000001010100000000000000000000000000000000000000000000110100000000001010000000000000011111000000000000111011111111111010101111111111101110111111111111011011111111111100001111111111111000111111111101001111111111111110110000000000000011111111111110000000000000000100101111111111111100000000000000001011111111111010000000000000000001111111111111001000000000000000101111111111100101111111111111111000000000000001010000000000001101000000000001000100000000000011000000000000010011000000000001001100000000000011011111111111101110000000000001100111111111111101111111111111111011000000000000011011111111111110101111111111110011111111111100101011111111110101011111111111110100111111111110010011111111111111111111111111101001111111111111101011111111111111100000000000000001000000000001010111111111111110001111111111111010000000000001011011111111111010000000000000001101000000000000100011111111111000011111111111111011111111111110101111111111111011110000000000001010111111111111100011111111111110000000000000001001111111111110100000000000000010110000000000011000111111111111000100000000000001011111111111010111000000000000100100000000000011001111111111111101111111111110101011111111111110000000000000000010000000000100000000000000001011001111111111100111111111111111000011111111111101011111111111100101111111111111001111111111111100000000000000000110000000000011111100000000000010101111111111011010000000000001011111111111111000101111111111101110000000000001011011111111111110111111111111100001000000000001111000000000000100001111111111111100000000000001000000000000000000001111111111101000000000000001000100000000000000011111111111111000000000000001100000000000000100010000000000000000111111111111001000000000000000000000000000000001000000000000001000000000000011110000000000000001111111111110111100000000000110000000000000011111111111111111111100000000000110111111111111111100000000000000100100000000000001001111111111101000000000000000101011111111111101101111111111111101111111111110101000000000000011111111111111111001111111111111001011111111111110011111111111110100111111111111100000000000000100001111111111110111111111111111111111111111111100111111111111110111000000000000010011111111111001011111111111110100111111111111100111111111111001111111111111111000111111111111001011111111111110001111111111111110000000000000101011111111111110001111111111110100000000000000011100000000000000110000000000010000111111111110110111111111111100110000000000000001000000000000101111111111111001000000000000001011000000000000001011111111111110110000000000000011111111111111011011111111111001001111111111111110111111111111111011111111111100011111111111111111111111111110111111111111111101010000000000100010111111111111101011111111111010110000000000010101111111111101101100000000000101100000000000011001000000000000100000000000000001001111111111101000000000000000011100000000000001111111111111111110000000000000000111111111111101111111111111101101111111111111111000000000000010100000000000001111111111111111111111111111111110111111111111111100000000000000001011111111111110001111111111111001111111111111010000000000000101000000000000000000111111111111010111111111111110011111111111110110111111111111101011111111111111000000000000000000111111111111111011111111111111101111111111111011000000000000001000000000000001001111111111110011000000000000100100000000001001001111111111110000111111111111110000000000000000001111111111111000111111111111101100000000000001011111111111110101000000000001010011111111111011101111111111101011111111111110111011111111111101000000000000000000111111111111001011111111111110100000000000000001000000000000000011111111111110011111111111110111000000000000000000000000000010011111111111111000111111111110001000000000000000101111111111101111000000000001000111111111111111111111111111111000000000000000000100000000000001101111111111110100000000000000000000000000000010001111111111110110000000000000101011111111111011001111111111111100000000000000110100000000000010001111111111111001000000000000010000000000000001001111111111100100000000000000000011111111111110101111111111010000000000000000110111111111111110010000000000000110000000000000000011111111111011001111111111111111111111111111111011111111111111010000000000000110000000000000001100000000000010111111111111111010000000000000001100000000000010111111111111110000000000000000000011111111111100111111111111111001111111111111101011111111111101110000000000000011111111111111011000000000000000100000000000000000111111111111011111111111111111100000000000000000000000000000001011111111111011001111111111110011000000000000000111111111111101101111111111111111000000000000001111111111111101010000000000000111111111111111000111111111111010100000000000010110111111111111010111111111111100100000000000010100111111111111011011111111111110110000000000101110000000000000110000000000000011011111111111110110000000000010010100000000000011011111111111110001111111111111100011111111111101111111111111101011000000000000000000000000000011100000000000001011000000000000100100000000000010011111111111111101111111111111110100000000000010010000000000001101000000000001110000000000000111110000000000010111111111111110111111111111111111011111111111010110000000000001010100000000000001110000000000001101111111111111000111111111110110001111111111100111000000000000010000000000000000011111111111110111000000000000011111111111111001010000000000001001000000000010000011111111111101010000000000001110000000000000001100000000000010111111111111101101000000000000101100000000000101001111111111100010111111111111100000000000000001100000000000011010000000000000001011111111111100110000000000011100111111111111110011111111111111000000000000001010000000000001010000000000000010110000000000010010000000000000000111111111110101001111111111111011111111111110110011111111111110001111111111110101000000000000111000000000000100001111111111101111111111111111010111111111111100101111111111101010000000000000001000000000000100100000000000001001000000000001000100000000000000111111111111110111111111111111111011111111110111111111111111011100000000000000000000000000000011100000000000001011111111111111010000000000000001101111111111101101000000000000111100000000000100011111111111101110000000000000001000000000000001001111111111101110111111111111110011111111111011110000000000000011000000000000000011111111111101100000000000000100111111111111001011111111111110010000000000001110000000000010110000000000000101011111111111011010000000000000010011111111111101110000000000001001000000000001111100000000000100010000000000000011000000000010100000000000000010100000000000000100111111111110111111111111111000101111111111111011111111111110000111111111111101001111111111101100111111111111111000000000000000110000000000001001111111111111011011111111111100001111111111110100111111111111110111111111111100111111111111101001000000000000111011111111111101111111111111110100111111111111100011111111111101101111111111110001000000000000111000000000000010011111111111111001000000000000011100000000000011010000000000001001000000000000000011111111111101011111111111111010111111111110110111111111111000111111111111010110000000000001011111111111111111100000000000000110000000000000010100000000000000111111111111111000000000000001011000000000000100010000000000000000111111111111101100000000000001100000000000000100111111111111111100000000000100101111111111110111111111111111101000000000000010011111111111011011000000000000101100000000000010000000000000101000111111111110010011111111111101110000000000100100111111111111011111111111111011101111111111111110000000000010110100000000000101100000000000010000111111111111101111111111111100110000000000000000000000000001100100000000000111111111111111110111111111111111101100000000000010101111111111110000000000000000011100000000000011000000000000000000111111111110100111111111111011000000000000000000000000000001101011111111111101011111111111101110000000000010000011111111111111011111111111101110000000000010000100000000000010101111111111101011111111111101111011111111111110000000000000001100111111111111010000000000000000010000000000011110000000000010001100000000000010101111111111110010111111111111011100000000000011000000000000010001111111111111111011111111111101001111111111110011111111111111001111111111111000111111111111100111111111111111100000000000000000000000000000011010000000000000100000000000000000010000000000001011111111111101110111111111111001011111111111111100000000000000000100000000000010011111111111101110000000000000000111111111111010100000000000000001000000000001000011111111111100001111111111101011000000000001110100000000000100101111111111111011000000000000000000000000000110000000000000001101000000000001010100000000000010101111111111101110000000000000000000000000000011110000000000101001111111111110111000000000000111001111111111110111111111111111011000000000000000111111111111011101000000000001010000000000000000000000000000000000000000000000001111111111110110001111111111110101000000000000000011111111111101110000000000000111000000000000001000000000000001101111111111011010000000000010000111111111111100011111111111101001000000000001001000000000000011011111111111101001111111111110110000000000000010101111111111110001111111111011110111111111111001001111111111111000111111111011101011111111111101100000000000101100000000000001111100000000000001100000000000010100000000000000000100000000000101100000000000000101111111111110001011111111111011011111111111110011000000000000110100000000001011011111111111110010000000000000010000000000001000110000000000000000000000000000101100000000000010101111111111101000111111111111111111111111111011100000000000000001111111111111111111111111111000110000000000011000000000000000011111111111111011110000000000000101111111111111111100000000000010110000000000000001111111111111001111111111111100111111111111111101000000000000000111111111111110010000000000011000000000000000101011111111111101001111111111111000000000000000011011111111111110000000000000000010111111111111110100000000000001000000000000000001111111111101111100000000000001111111111111110000111111111110001000000000000000011111111111101001111111111101010111111111111011101111111111111111000000000000001011111111110111110000000000001001000000000000000000000000000001000000000000101000000000000001001100000000000111110000000001010000000000000000111111111111111011111111111111110011111111111111000000000000000001000000000000011110111111111111011100000000000101010000000000110001111111111110000111111111110111111111111111100111111111111101001000000000000000000000000000000000111111111101100100000000000010110000000000000111000000000001000011111111111111001111111111011101111111111111011011111111110111101111111111100110111111111110001011111111111101101111111111101001000000000000000000000000000000001111111111110101111111111110110011111111111110101111111111101110111111111111011111111111111110111111111111110011111111111111000000000000000000001111111111100110000000000000001011111111111011001111111111000101111111111110110011111111111011101111111111001001000000000010110000000000000100011111111111011001111111111111101100000000000000001111111111111101111111111111010100000000000000101111111111111010000000000001100100000000000100011111111111111101111111111111000100000000000000100000000000000001000000000000110100000000000110011111111111111110000000000001011000000000000101001111111111111101111111111111110111111111111111111111111111111100111111111111111111111111111100001111111111101011111111111111111011111111111100001111111111011101000000000000111000000000000010011111111111101100111111111111010011111111111110001111111111110011111111111110011011111111111010010000000000000010111111111110111000000000000110100000000000001111111111111101101100000000000110110000000000001010111111111110110000000000000000111111111111111001000000000010000100000000001011000000000000010010000000000010011000000000000110101111111111001001000000000000000111111111111110010000000000100010000000000000100100000000000001100000000000100011111111111111101000000000000001100000000000001100111111111111110111111111110100101111111111101111111111111110101111111111110101110000000000000001000000000001010100000000000000100000000000001010000000000000101111111111110111011111111111010100000000000001011111111111111110011111111111110010000000000001110011111111111111101111111111100110111111111111000000000000000000110000000000010110000000000000101011111111111010000000000000010101000000000000000000000000000110100000000000000100111111111111101100000000000010101111111111111101111111111111001100000000000001000000000000001110111111111111101000000000000011110000000000000110000000000000001100000000000100100000000000001001000000000000100100000000000000111111111111111001111111111101111011111111110101101111111111100011111111111111101011111111111011000000000000000111111111111111000011111111111111100000000000000001000000000001001000000000001000100000000000010100000000000001010111111111111100000000000000000000000000000000000011111111110111001111111111101110000000000001101000000000000101110000000000000100111111111110101011111111101110111111111111001010000000000001010111111111111101100000000000011100000000000001001000000000001010110000000000010100111111111111000011111111111110101111111111110110000000000000001100000000000101100000000000000000111111111111011111111111111010100000000000000111000000000000000011111111111110110000000000100111111111111111111100000000000010110000000000100000111111111111000011111111111111101111111111111011000000000000001100000000000010101111111111111010000000000010010011111111111110110000000000010110111111111101110111111111111010011111111111110101000000000001010011111111111110100000000000011101111111111111101111111111111100001111111111101011111111111101111011111111111001101111111111111011111111111111110000000000000111110000000000100111000000000000011000000000000000000000000000001011111111111111011011111111111011010000000000000000000000000001000100000000000001100000000000000001000000000000011000000000000010000000000000001011111111111111110011111111110101101111111111100000111111111110011100000000000011100000000000011101000000000000101100000000000010010000000000100000000000000010101100000000000110110000000000000010111111111110101011111111111000101111111111111111111111111111111000000000000000000000000000010111000000000001000000000000000000000000000000001100111111111110111011111111111111011111111111111011111111111111000000000000000010010000000000110101111111111110100111111111111100110000000000000000111111111011110011111111111001000000000000010110111111111110111111111111111111110000000000111010000000000001010000000000000011010000000000010100000000000001110011111111111000101111111111110100000000000000001111111111111100011111111111110110111111111111111111111111111101011111111111101001111111111101110011111111111011101111111111110110000000000000000100000000000011110000000000001000000000000001000100000000000000100000000000000100000000000000000100000000000000001111111111010110111111111111011000000000000010110000000000001001000000000001111100000000000010000000000000010011000000000001101011111111111111101111111111010111000000000000000000000000000001000000000000011110000000000001000111111111111101011111111111101110000000000011000011111111110011111111111111100001000000000000001011111111111101011111111111011101000000000000111011111111111011111111111111100011111111111111000111111111110111011111111111100000111111111111000111111111111011011111111111101110000000000000111000000000000011111111111111111100;
endcase
end
endmodule



module lut_weights_6(sbyte,addr);
input [3:0] addr;
output reg [82943:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0110: sbyte = 82944'b111111111111011111111111110110011111111111100111111111111110110011111111111100000000000000001001000000000000111111111111111111111111111111110000000000000000010011111111111100110000000000000101000000000000100111111111111101001111111111110001111111111111000111111111111110000000000000001010111111111111100011111111111110111111111111110010111111111111001100000000000010010000000000000111000000000000010100000000000000100000000000011010111111111111111000000000000000000000000000001001000000000000111000000000000100001111111111111100000000000000010111111111110111100000000000000000000000000000010000000000000011000000000000000101111111111111011011111111111110101111111111101101111111111111100111111111111110101111111111110111000000000000001111111111111110001111111111110111000000000000111111111111111110010000000000000111000000000000000000000000000011011111111111101000111111111110110111111111110111101111111111110101111111111110100111111111111100111111111111011100000000000010001000000000001001011111111111111010111111111111111111111111111111110000000000010100111111111111010000000000000100111111111111110000000000000000011011111111111110011111111111100000000000000000111000000000000000001111111111111111000000000000001000000000000100110000000000010010111111111110111000000000000110000000000000100111111111111111010111111111111101010000000000000100000000000000110111111111111110001111111111111111111111111111101000000000000001011111111111111111111111111111100111111111111110011111111111110000111111111111001111111111111010101111111111100000000000000000101011111111111011111111111111110101111111111111110011111111111011011111111111110101111111111111011011111111111110101111111111110101111111111111111100000000000010101111111111111100000000000001000000000000000100100000000000001001000000000000100111111111111110110000000000000111000000000010011000000000000101000000000000001010000000000010001000000000001001100000000000001101111111111111011111111111111101101111111111111111111111111111101111111111111110001111111111101111000000000000111000000000000011010000000000010110111111111111100000000000000001110000000000000001111111111111010100000000000001000000000000001101111111111111011000000000000011010000000000010000000000000001111011111111111110011111111111110011111111111111001000000000000100010000000000010010000000000000000011111111111100011111111111101001111111111111010000000000001000001111111111111011000000000000101011111111111111010000000000000011111111111101111111111111111000101111111111110010111111111111111111111111111110101111111111101110000000000000001100000000000111010000000000010100000000000000010000000000000001100000000000000000000000000001011011111111111011000000000000000111000000000100000100000000000110100000000000010100000000000000000011111111111011001111111111100111111111111111100111111111111011101111111111101000111111111111100011111111111110110000000000000011000000000000001011111111111101101111111111111001111111111111100100000000000001111111111111111111111111111111011100000000000001011111111111110000000000000001010111111111111111110000000000000001111111111111010111111111111001010000000000001011111111111110011011111111111011111111111111110010111111111110111111111111111010011111111111111000111111111111011011111111111111101111111111110001000000000001000111111111111101011111111111111111111111111111110000000000000001011111111111111110111111111111100111111111111011111111111111111011111111111111100011111111111111011111111111110110000000000001011000000000000100010000000000101000111111111110111111111111111100110000000000000000111111111110111011111111111110010000000000010111000000000001011100000000000011111111111111111101111111111111001100000000000010111111111111111110000000000001100011111111111110101111111111111110111111111111011111111111110111010000000000000100111111111101000011111111110111001111111111101111111111111110010111111111111010100000000000000010000000000011010100000000000011100000000000000100000000000010111111111111111111011111111111111100000000000000100111111111111110000000000000000011111111111111011000000000000010101111111111110000000000000001001000000000000000101111111111011101000000000000100111111111111010101111111111010100111111111111000111111111111101100000000000001110000000000000110011111111111111011111111111111010111111111111110011111111111110001111111111110111000000000000000100000000001000100000000000101011000000000001101100000000001011000000000000010100000000000000111111111111111110101111111111011101000000000000101000000000000100101111111111011011000000000001111100000000000100001111111111111010000000000001111100000000000000100000000000011101111111111111111011111111111100111111111111110011111111111110000111111111111010011111111111100100111111111110010000000000000000111111111111111001111111111111100100000000000010111111111111111000000000000000011100000000000101010000000000010010000000000001010111111111111111100000000000000101111111111101010011111111110101101111111111010100000000000000010011111111111100011111111111000111000000000001111100000000000001011111111111101110111111111111111111111111110100111111111111001011000000000000101111111111111111001111111111111101000000000000001111111111111011110000000000000100000000000001001011111111111111111111111111111101111111111110101000000000000000110000000000000100111111111111010000000000000000011111111111111111000000000000000000000000000010111111111111110111111111111110111111111111110111011111111111101111000000000000111111111111111001011111111111110011111111111110111100000000000001010000000000001010111111111111111011111111111111010000000000000111000000000000001100000000000010000000000000010001000000000000110011111111111000001111111111101100000000000000000100000000000001000000000000010011111111111110010100000000001000000000000000101010111111111101001111111111110101111111111111010011000000000000010000000000000010010000000000001101000000000001100100000000001000000000000000101111111111111110000011111111111010110000000000010101000000000011001000000000000110101111111111110100000000000011101000000000000100101111111111111111000000000001101011111111111011010000000000101010000000000010101111111111111100111111111111111111111111111101101111111111111110010000000000010100111111111110100011111111111011001111111111110111111111111110011011111111111000011111111111111000000000000001001000000000000101010000000000101001000000000001100100000000000010111111111111111101000000000001110000000000000100101111111111110001000000000000101100000000000000011111111111111000111111111111111111111111111111010000000000000001000000000001100000000000000000101111111111111111000000000001100111111111111010100000000000000000111111111101101011111111111010010000000000000000000000000000110111111111111010001111111111011111000000000001010111111111111010011111111111011100111111111110111100000000000101110000000000010010111111111111110000000000001000000000000000100110111111111110100011111111111111100000000000100001000000000010010100000000010000000000000000100010111111111100010000000000000000000000000000110100111111111110001111111111111011110000000000011001111111111111110111111111111011100000000000001100111111111111101000000000000001010000000000000110000000000000100000000000000100101111111111110111111111111111100000000000000010111111111111101000111111111101001111111111111000101111111111111110111111111110101011111111111001001111111111110000000000000001010000000000000100111111111111101110000000000011001011111111111010111111111111101101000000000010010011111111111111100000000000001100000000000000101111111111111001111111111111010101000000000001111000000000000001111111111111100010111111111111111100000000000101001111111111111000111111111111110100000000000001101111111111101011111111111110001100000000000001110000000000000000111111111101101011111111111011101111111111110000111111111111100011111111111100110000000000011100000000000001100111111111111101100000000000000001000000000000100111111111111101101111111111101011111111111101001100000000000100000000000000101001111111111101100011111111110000110000000000000101000000000000010011111111111111100000000000000111111111111111010111111111111100001111111111011100111111111111011100000000000000001111111111111010000000000000010000000000000000001111111111101011111111111111100111111111111111000000000000001011111111111111001000000000000001011111111111111000000000000001011011111111111100110000000000001010111111111111011111111111101101001111111111001011111111111111111100000000000000101111111111111010111111111111100000000000000100001111111111110101111111111110101111111111111101111111111111111111000000000000100000000000000111100000000000000100000000000000101111111111111010101111111111011100111111111110111111111111111001101111111111111111111111111111000111111111111010111111111111011111000000000001101111111111111101111111111111100001000000000000110011111111111010011111111111010100000000000000101111111111111111101111111111111010000000000000000000000000000001111111111111111100111111111110100011111111111000101111111111111110111111111111000100000000000000101111111111111100111111111110111000000000000000111111111111110100000000000001101000000000001010000000000000011000111111111101111100000000000000110000000000001100111111111111000011111111111010010000000000010100000000000001111100000000001001010000000000101100111111111111100100000000000000110000000000001100111111111110100011111111110110001111111111110001111111111110110000000000000100001111111111110010000000000000110011111111111011010000000000001111000000000000011100000000000100000000000000100000000000000001100000000000000000011111111111111001000000000000010111111111111101111111111111111001000000000000000000000000000000110000000000000001000000000010100100000000000111000000000000000011000000000000000000000000000000100000000000001000000000000000000011111111111100001111111111110001111111111110000011111111111111101111111111111110000000000010000100000000000000011111111111100111000000000001100000000000000010111111111111101111000000000010000100000000000000101111111111011110000000000000000111111111111011010000000000000111111111111110100100000000000100100000000000011100000000000000010011111111111010011111111111100101000000000010010000000000000001100000000000000110000000000010011111111111111101010000000000000111000000000011000000000000011000000000000000010110000000000000101000000000000000100000000000001010111111111111000011111111111111010000000000011110000000000010010000000000000110100000000000011111111111111110101011111111111101001111111111111101111111111110111011111111111110011111111111110100111111111111111011111111111011000000000000000000111111111111110011111111111110011111111111111101111111111111100000000000000010110000000000000011000000000000010100000000000110111111111111111011000000000000111011111111110110001111111111011011111111111111101111111111111110010000000000001001000000000001100100000000001000100000000000100111000000000010100000000000001101000000000000011000000000000001110100000000000000001111111111100111000000000000001000000000000010000000000000100000000000000000001111111111111101110000000000001010000000000000011100000000000010111111111111111111000000000000000111111111111111001111111111111011000000000000001000000000000001000000000000001110111111111111101100000000000001111111111111101110000000000000000011111111111101011111111111111011111111111111000100000000000000001111111111110110111111111110101111111111111011110000000000000000111111111110100011111111111110011111111111111100000000000000001100000000000110000000000000010100111111111111011111111111111101111111111111101010111111111111100000000000000001001111111111110100111111111111011111111111111111101111111111101110000000000001010111111111111010111111111111111000000000000000001000000000000011001111111111110101111111111111001000000000000101001111111111101011111111111111011000000000000001100000000000010010000000000010001000000000000101100000000000011001111111111111110100000000000100100000000000110000000000000001101000000000000101101111111111111101111111111111100000000000000010010000000000011010111111111111010011111111110111011111111111110111111111111111010011111111111010110000000000000111000000000000101000000000000000001111111111101110000000000000111111111111111111001111111111100010000000000000111100000000000001011111111111010001000000000000011111111111111111100000000000001111111111111110110111111111111101100000000000010001111111111101100000000000000010010000000000010010000000000010000111111111110111011111111111101110000000000001000111111111111100011111111111100110111111111111100011111111111010111111111111110011000000000001001100000000000000000000000000000111000000000010001000000000000100000000000000000000000000000000010100000000000010011111111111110101111111111110001111111111110101001111111111101011111111111111110111111111111110000000000000010101111111111111110000000000000010100000000000110011111111111110110100000000000001000000000000000001000000000000000011111111111010110000000000001000111111111111000011111111111010100000000000000100000000000010010100000000000011001111111111101010000000000000111111111111111101101111111111011110111111111111010111111111111100001111111111011000000000000001000100000000000001100000000000001000111111111101101011111111111000011111111111001101111111111110101111111111111000001111111111110000111111111110111000000000000110101111111111101111000000000001001111111111111101110000000000011001000000000000001011111111111101110000000000001000000000000000000011111111111100101111111111101011000000000000111000000000000010111111111111110001111111111111011000000000000011011111111111111001111111111111001011111111111100001111111111100001000000000000010011111111110111011111111111101110111111111111001011111111111110010000000000000010000000000000011100000000000000110000000000011110111111111111001100000000000001010000000000001100111111111111110100000000000011000000000000000000000000000011001000000000001110010000000000110010000000000001000100000000000010011111111111111110000000000000000011111111111010011111111111110100000000000000100000000000000001100000000000001110000000000000011011111111111111010000000000000111111111111111100100000000000100100000000000000111111111111111100111111111110111111111111111110000111111111111111011111111111001011111111111111010111111111111000100000000000000000000000000001111000000000011000111111111111100011111111111111011000000000010000000000000000010000000000000011100000000000001011100000000000100110000000000001111111111111111100100000000000010011111111111110010000000000010011100000000000010110000000000001010000000000000001000000000000000011111111111111110000000000000010011111111111101011111111111110101111111111111101111111111111010100000000000011010111111111111100111111111111011001111111111101110111111111111010100000000000010111111111111011000000000000001011000000000001000101111111111110011111111111111100000000000000001101111111111110111111111111111000111111111111010011111111111110111111111111111101100000000000001000000000000001000000000000000011111111111111101100000000000010001000000000001110100000000000100000000000000000000000000000010010000000000000000001111111111110011111111111101100111111111111011111111111111101100000000000000011000000000000000000000000000000000111111111111110000000000000000011111111111101100111111111110111011111111111110100000000000000010000000000000011000000000001010000000000000100001000000000000011100000000001010110000000000001111000000000000010100000000000011100000000000001000000000000000001100000000001000000000000000011101000000000001011000000000000110100000000000001011000000000000110011111111111100011111111111111111111111111110100111111111110000111111111111010001000000000001100111111111111110011111111111100100000000000000000111111111111110011111111111110100111111111110010011111111111000011111111111101000111111111111100000000000000110110000000000000100111111111111100000000000000010010000000000001011111111111110111011111111110111101111111111110100111111111111101011111111111101111111111111111101000000000000110011111111111010110000000000011001111111111111001111111111111011101111111111100110111111111111101011111111111100001111111111111111000000000000111100000000000010110000000000010000000000000000000000000000000110110000000000110011111111111111011011111111110111111111111111101010111111111100000111111111110110100000000000001011111111111110101011111111111011000000000000000000111111111111101111111111111100111111111111111000000000000001111000000000000011011111111111110101000000000001100011111111111000111111111111100101000000000010000100000000000000101111111111111100000000000010000100000000000000001111111111111100111111111110100000000000000000000000000000010000111111111111111111111111111111010000000000001111111111111110110011111111111100001111111111101011000000000001111011111111111100110000000000101000000000000000001100000000000100100000000000001010000000000000111111111111111111010000000000001101000000000010101011111111111100111111111111010110111111111110100011111111111110100000000000010111000000000001100100000000000000100000000000000101000000000000110111111111111110001111111111110101000000000001001000000000000110001111111111111000000000000000101100000000000100011111111111101100111111111101100011111111111001011111111111101011111111111101101011111111110111111111111111110100111111111110010011111111111001111111111111111100111111111111111000000000000001001111111111101000111111111111001000000000000110010000000000010110111111111111110100000000001010000000000000010000111111111111010000000000000011000000000000000110000000000000100000000000000010110000000000001110111111111111110000000000000000000000000000000101000000000001000000000000000101000000000000011001111111111111011000000000000010000000000000010000000000000000111000000000001000110000000000100010111111111111100011111111111111001111111111110011111111111110011100000000000011011111111111111110111111111110010111111111111110101111111111101100111111111101110011111111111111110000000000000110000000000000000011111111111000001111111111010111111111111110001011111111111011111111111111011100111111111110111000000000000110100000000000000100111111111110101000000000000000110000000000001111111111111011011011111111101010101111111110100110000000000010100011111111111110111111111111110010000000000000000100000000001001011111111111110100000000000001101111111111111110000000000000100000111111111111110011111111111111110000000000001011111111111111111100000000000011000000000001001010111111111110001111111111111101111111111111100111000000000000011111111111111011100000000000010100000000000001010111111111111101010000000000001011000000000001110100000000000100000000000000001010111111111111101000000000000001001111111111110001000000000000000111111111111010111111111111111011111111111110111100000000000001001111111111110101111111111111010000000000000000000000000001001100000000000001100000000000000011110000000000011001000000000001010111111111110110101111111111010000111111111111111011111111111101011111111111111010111111111111100111111111111010011111111111111010111111111111010100000000000001001111111111101100000000000000100000000000000000001111111111100110111111111111011011111111111110001111111111101011111111111110100011111111111011101111111111100110000000000000000011111111111110010000000000010100111111111111011111111111111101111111111111101100000000000000011011111111111001011111111111100101111111111110100111111111111100001111111111100000111111111111001011111111111110101111111111111101000000000001010000000000000111000000000000100011000000000010000000000000001000100000000000001100000000000000010011111111111111001111111111110100000000000001101011111111111011101111111111100000111111111111010100000000000011100000000000110111111111111111010000000000000101000000000000011010000000000001111000000000000100110000000000100001000000000000010100000000000101010000000000001000111111111111110111111111111010001111111111111101111111111110100111111111111111001111111111101011000000000000010100000000000000111111111111101011111111111110110000000000000000101111111111010011111111111111000111111111111011011111111111110111000000000001100011111111111101001111111111101100000000000000111100000000000011001111111111011000111111111111010011111111111011110000000000010000111111111111100100000000000001001111111111111111000000000000000000000000000000001111111111110001111111111111011000000000000001110000000000000000000000000000111000000000000100110000000000001010000000000001110100000000000000001111111111111100000000000000100111111111111110010000000000000011111111111111101011111111111100001111111111100101111111111110010011111111111111111111111111110010000000000001011000000000010000110000000000000100000000000000110111111111111101111111111111110111111111111111111000000000000001111111111111111001111111111111101011111111111101001111111111110001000000000000001011111111111010110000000000000011000000000001011111111111111110011111111111110001000000000000110000000000000000001111111111110000000000000000001011111111111101010000000000000101000000000000000011111111111111001111111111111101111111111111101000000000000011011111111111111100111111111111100111111111111101011111111111111011111111111111101011111111111110111111111111111110000000000000100111111111111011110000000000001111111111111111100100000000000000111111111111100011111111111111000111111111111111110000000000000000000000000000001000000000000000000000000000001000111111111110111000000000000011011111111111111101111111111111100100000000000001000000000000001010000000000001100100000000001000011111111111111111000000000001010000000000000111010000000000010110000000000000100011111111111101011111111111111000111111111110010111111111111101010000000000000111111111111100110000000000000000000000000000000110111111111110111100000000000100001111111111100101111111111111001011111111110111001111111111111100111111111110001000000000000000001111111111111101000000000001000111111111111001111111111111101010111111111111000111111111110110011111111110111111111111111111011111111111111001101111111111100011000000000001001000000000000110010000000000000001000000000011010100000000000110000000000000011000000000000001000000000000000101100000000000000001111111111111111011111111111111110000000000000011000000000000110111111111111101110000000000000000111111111110010000000000000001001111111111011110111111111111010111111111111101011111111111110000111111111110010011111111111110101111111111000101000000000001010100000000000110100000000000000011111111111111110111111111111110101111111111111110000000000000110100000000000011111111111111101101111111111101111011111111111101100000000000001101111111111111011100000000000000110000000000000100000000000000000100000000001000110000000000111010000000000000110000000000000100000000000000000111000000000000000000000000000010000000000000001001000000000000010000000000000110010000000000010101000000000000110011111111111110011111111111110110000000000001100011111111111110001111111111101001000000000001110000000000000101110000000000010111000000000001100100000000001100100000000000001101111111111111010000000000000000001111111111101101111111111101001011111111111110011111111111110010000000000000111000000000000011010000000000001011000000000001010100000000000010001111111111101100000000000000111011111111111010011111111111010100000000000000101011111111111001111111111111101100111111111111110111111111111010011111111111011100111111111101111111111111111010111111111111001010111111111111100011111111111110001111111111111000111111111110010000000000000100000000000000100001111111111111011100000000000001000000000000100011000000000011010000000000000110111111111111111100000000000001101000000000000101100000000000000101000000000001001111111111111101101111111111111001000000000000101100000000000011001111111111110001000000000000010011111111111101010000000000000010000000000010111011111111111110101111111111111100111111111110101111111111111111111111111111111110111111111111000100000000000010001111111111110001000000000000010100000000000100011111111111100011000000000000101111111111111110101111111111111000000000000010110000000000000111111111111111110110000000000011011000000000000111111111111111101110111111111111010100000000000100001111111111111111000000000000111000000000000000100000000000100000000000000001001011111111111111111111111111101000111111111101011011111111111000101111111111111010111111111101010111111111110110010000000000000000000000000000001111111111111010101111111111111111000000000000100011111111111111011111111111110000000000000000101100000000000001001111111111111001000000000000000000000000000101001111111111110001111111111110101111111111111111010000000000001111111111111110000100000000000001110000000000101000000000000000100000000000000001100000000000001100000000000001011111111111111110101111111111101101111111111110111000000000000000011111111111111110111111111111111111111111111101100000000000001010111111111111100100000000000101010000000000000001000000000000011000000000000001110000000000001000111111111111001111111111111100001111111111101010000000000000101100000000000000010000000000000000111111111111111100000000000000001111111111111000000000000000000011111111111010000000000000001000000000000001010111111111111011011111111111100000000000000010011000000000000100011111111111110000000000000001100111111111111100110000000000100001111111111111111111111111111110101111111111111000111111111111001000000000000001011111111111111111000000000001011100000000000011101111111111110101111111111111111011111111111010010000000000001101111111111111000000000000000010100000000000011110000000000000001000000000000000001111111111100111111111111110110011111111111111010000000000001000000000000000001100000000000001000000000000001001000000000000001000000000000000100000000000000101111111111111011000000000000011100000000000000001111111111111110100000000000001110000000000010010000000000000000000000000000000010000000000001000111111111111010000000000000001110000000000010000000000000000111000000000000011110000000000011011111111111111010111111111111110100000000000000000000000000000011000000000000010010000000000001011000000000000011000000000000000100000000000000100111111111111111111111111111100110000000000001010000000000000010000000000001010000000000000111010111111111111111100000000000100110000000000011000000000000000111011111111111010000000000000001111111111111111100111111111111010001111111111100011111111111110001011111111111001111111111111100101000000000000110011111111111101110000000000001101111111111111111000000000000110000000000000000011111111111111111111111111111100111111111111110111000000000001000100000000000000001111111111111100000000000001001000000000000001100000000000010101111111111110111100000000000000011111111111111000111111111110000111111111111110010000000000000000111111111110111111111111111000001111111111111010111111111111111111111111111101011111111111101010000000000000101111111111111110011111111111111101000000000001010011111111111001101111111111101000000000000001001111111111111110101111111111110111111111111110011011111111111100101111111111111110111111111111011111111111111000010000000000001110111111111110111100000000000011110000000000101000111111111111111111111111111100000000000000000101000000000000100000000000000001001111111111110011000000000000010100000000000100010000000000010001000000000000010111111111111111111111111111111001111111111101001100000000000101100000000000011110111111111101101011111111111111000000000000001100111111111111111011111111111111110000000000100010000000000001001011111111111110100000000000000011000000000000101111111111111111101111111111110100000000000000011011111111111010011111111111110110000000000000010011111111111111100000000000010111000000000000100100000000000001110000000000001110000000000001001000000000000000101111111111110111111111111111110000000000000101110000000000101110000000000000011100000000000110110000000000000101000000000000011100000000001010000000000000000110111111111111111011111111110111110000000000000000000000000001010111111111111110000000000000000110111111111110101100000000000010111111111111111110000000000000101000000000000001011111111111011110000000000000100000000000000000001111111111010011111111111111111111111111111100011111111111011011111111111101110100000000000100010000000000000101111111111111010100000000000011000000000000000011111111111101001011111111110111001111111111110110111111111111110111111111111100110000000000001000111111111111101100000000000101010000000000000100000000000000100100000000000100010000000000000100000000000001001000000000000000101111111111111001111111111111011011111111111100101111111111100111111111111110000011111111111001011111111111100010000000000000001011111111111100010000000000100000111111111110001111111111110000011111111111011000111111111110011011111111110111010000000000010001000000000010011000000000000010010000000000000001111111111110100011111111111011010000000000000001000000000000000111111111111010001111111111101100111111111110011011111111111100101111111111110010111111111111100011111111111010101111111111101011000000000001001000000000000011001111111111110000111111111111110100000000000010000000000000010101000000000000000111111111111111101111111111101101000000000000011100000000000000110000000000000001111111111110000011111111111111010000000000000111000000000001001011111111111110101111111111111000000000000000101100000000001101000000000000011110000000000000111100000000000111010000000000000011000000000001000100000000000000100000000000001111000000000000111100000000001011010000000000111100111111111111011000000000000001111111111111111110000000000000000111111111111010001111111111010000000000000010100011111111111000011111111111001111111111111111010100000000000101100000000000000000000000000000000000000000001000100000000000000110000000000001110000000000001101110000000000001111000000000000101100000000001000110000000000010011000000000001001000000000000011000000000000000000000000000000101000000000000001011111111111101100000000000001000011111111111110111111111111101001111111111111010011111111111011001111111111011100000000000000101011111111111011011111111111100110000000000000101100000000000000011111111111110001111111111111001100000000000001101111111111110001000000000000010100000000001011001111111111111001000000000001101111111111111111110000000000000101000000000001010100000000000010110000000000010001000000000001011000000000001010110000000000111110111111111111100111111111110101011111111111011110111111111111001000000000000011001111111111110001111111111111101011111111111111011111111111000110000000000000111100000000000101010000000000101001111111111101111111111111111111000000000000000100111111111111101011111111111111110000000000000010000000000001000100000000000011000000000000000100000000000000111000000000000010100000000000011010000000000000101100000000000101010000000000001001000000000000111100000000001001101111111111011010000000000000111000000000000011111111111111111001000000000000100011111111111101001111111111001100111111111111111011111111111100011111111111110100111111111111010100000000000000111111111111110110000000000000110100000000001100100000000000001001000000000001100111111111110111111111111111100000000000000000011011111111111111101111111111011111000000000000000011111111110111001111111111010010000000000010000100000000000100101111111111110101111111111111000000000000000001001111111111110010000000000001001000000000000000011111111111110000000000000000010111111111111100100000000000001110000000000001000000000000000000001111111111110111000000000000010111111111111111011111111111111111000000000000010000000000000001000000000000001101000000000010001111111111111111110000000000000011111111111111010000000000000100110000000000000001000000000000100111111111111111001111111111111111000000000000110100000000000010110000000000000001111111111110010000000000000000010000000000100010000000000001011111111111111101011111111111100011000000000000101100000000000011000000000000000100000000000000100100000000000000010000000000000000000000000000001100000000000000001111111111110011000000000000011011111111111011101111111111111010000000000000000011111111111111101111111111111011000000000001101100000000000000001111111111010110000000000001011000000000000110000000000000100101111111111111111111111111111110010000000000001010000000000001001111111111111011011111111111111111111111111111010111111111111110000000000000011000111111111110000100000000000000010000000000001011000000000001111100000000001000110000000000011001000000000000011011111111111010111111111111110111000000000000010111111111111111000000000000000000000000000000000011111111111101000000000000001000000000000010000011111111111111110000000000001001000000000000000000000000000011101111111111110001000000000001000111111111111010111111111111010111111111111110111011111111110111011111111111100110000000000000000011111111111111010000000000010100000000000001110011111111111000111111111111101101000000000000011011111111111011100000000000000111111111111111110000000000000001111111111111101000000000000000000000000000000010110000000000001011000000000001011011111111111111110000000000010010111111111111011011111111111011100000000000000011111111111111101011111111111010011111111111110110111111111111010111111111111111111111111111011110111111111110111111111111111001001111111111100000000000000001100000000000001001010000000000011111111111111111111000000000000101000000000000011100000000000000100111111111111100110000000000000110000000000000010011111111111000101111111111001011111111111111100100000000000010001111111111110110000000000010000100000000001000010000000000001001000000000000001000000000000001011111111111110000000000000000110011111111110100001111111111100000000000000001101000000000000000001111111111111000000000000000000111111111111111011111111111111101000000000001000000000000000010010000000000010100111111111101110011111111111101011111111111011000111111111111100011111111111111001111111111111110000000000000110100000000001000100000000000001100111111111110011111111111111110010000000000100100000000000001011000000000000001011111111111010111000000000000110000000000000000111111111111100110000000000000010000000000001001100000000000001011000000000001110111111111111111001111111111111110000000000000001100000000000001100000000000000010111111111111010011111111111101011111111111111011000000000000011111111111111101100000000000000000000000000000111111111111111110111111111111101101000000000000111000000000000011100000000000000101000000000001010011111111111101111111111111101001000000000000010100000000000010000000000000000000000000000001111011111111111111000000000000000110000000000000000100000000000100010000000000010011000000000000110000000000000110000000000000000110000000000001100000000000000010100000000000000100111111111110110011111111111010001111111111010010111111111110101011111111110101111111111111111010111111111110101000000000000000000000000000010100111111111111000100000000000010111111111111110000000000000001001100000000000110010000000000010101000000000000101100000000000010100000000000000110111111111110000100000000000001010000000000001000111111111101110111111111111110011111111111111001111111111110101111111111111011110000000000010000000000000001010000000000001000111111111111110010111111111110011000000000000001000000000000001000111111111110111011111111111110010000000000001011000000000000001100000000000010100000000000000001000000000000001000000000000100101111111111110100000000000000000100000000000010000000000000001110111111111110110000000000000010011111111111111101111111111111111000000000000011110000000000010011111111111110111011111111111011100000000000000000111111111110000011111111111001011111111111100100111111111101100011111111111001110000000000000000111111111111100111111111111111011111111111100000111111111111011100000000000111100000000000011111000000000001011000000000000001001111111111110001000000000000111011111111111111100000000000000111111111111110010011111111111011110000000000000101111111111100011011111111111111010000000000001111111111111110010111111111111100101111111111111101111111111111101011111111111011111111111111111011111111111111011000000000000001010000000000000101000000000000111100000000000000100000000000000110000000000000000111111111110111001111111111011010000000000000011011111111111110111111111111100101111111111111101011111111111101101111111111111010000000000000111111111111111101000000000000000010000000000000000000000000000000001111111111101001111111111111000111111111111011011111111111110101000000000010000100000000001001110000000000101011111111111111100000000000000100110000000000000111000000000000000011111111111101001111111111110000000000000011010000000000000111010000000000100110000000000001101100000000000000000000000000011011000000000010010000000000000110000000000000010011000000000000000000000000000011010000000000000110000000000000111100000000000000010000000000001111111111111111010100000000000101010000000000000011000000000000010000000000001000110000000000011100111111111110111011111111111011011111111111110111111111111110000111111111110110100000000000000011111111111110010011111111111100001111111111111111111111111110110100000000000010000000000000001001000000000000000011111111111110100000000000001100000000000000000011111111111111111111111111111100000000000000110000000000000100010000000000001011000000000010100000000000001000111111111111111000111111111111111000000000000001110000000000010010111111111111010000000000000001100000000000100001111111111111011111111111111001001111111111110100111111111111101111111111111111101111111111111101111111111101101111111111110111101111111111100101111111111100100111111111111000110000000000000000000000000000011100000000000000100000000000001111000000000000100000000000000000000000000000010100000000000001011111111111111110100000000000001001111111111100100100000000000001000000000000011110111111111100011000000000000000000000000000101101111111111110100000000000000010110000000000001100111111111110010111111111110101001111111111110011000000000000011011111111111101011111111111110010000000000001100111111111111111111111111111110111000000000000111000000000000010010000000001001001111111111111010100000000000011000000000000000110000000000000000111111111111101011111111111110110111111111111001011111111111011101111111111110101000000000000001100000000000011011111111111101101111111111111110100000000000101111111111111101011111111111111001100000000000001011111111111110100111111111111110000000000000010011111111111111011111111111111011100000000000011100000000000000010000000000001010000000000000101100000000000000100000000000001111111111111111101111111111111011001111111111111101011111111110011011111111111001001111111111111011100000000000001011111111111101110000000000001010100000000000011110000000000001001000000000100010100000000000111000000000000000000000000000000001111111111111011111111111111011011000000000000100111111111111111111111111111101110000000000001111100000000000111011111111111101010000000000000111100000000000011100000000000000101111111111111111111111111111100000000000000010100111111111111010011111111110110001111111111110101111111111110010011111111111111000000000000101000111111111101101011111111111011001111111111100100111111111110111111111111111010101111111111111100000000000001001111111111111101111111111111101001111111111101101011111111111010111111111111011110000000000001011111111111111101101111111111111001000000000001010000000000000011111111111111100110000000000000010011111111111110101111111111100110000000000000110111111111111000011111111111010000000000000000111100000000000011001111111111111100000000000001101011111111111110010000000000001000111111111111001100000000000000000000000000001000111111111111000111111111110110011111111111101011111111111111001011111111111100010000000000000001000000000001001000000000001000000000000000011110111111111111101000000000000000001111111111110010111111111111001111111111111101010000000000001011000000000000100111111111111111110000000000011100111111111111011011111111111100101111111111111000111111111111111111111111111111111111111111110010111111111111010000000000000001001111111111110110111111111110001011111111111010101111111111100110000000000000101000000000000111001111111111110001000000000001000000000000001000000000000000000000111111111111111111111111111101101111111111110001111111111111100011111111111011001111111111110101000000000001000011111111111110101111111111101110000000000000100011111111111101011111111111111010111111111111001000000000000010100000000000010010111111111110110000000000000100000000000000100000111111111110111011111111111100001111111111100000000000000000001011111111111111000000000000010000111111111111010100000000000101000000000000010011111111111110100100000000000000000000000000010100111111111111110100000000000100101111111111100111111111111101101100000000000000110000000000000011111111111111100000000000001000100000000000010110000000000000101111111111111100011111111111010100000000000000110100000000000001101111111111011110111111111111100100000000000010110000000000000100000000000000011011111111111010110000000000000001111111111111001011111111111000111111111111101011111111111111111100000000000101000000000000000011111111111111101000000000000100100000000000010011111111111111100111111111111101110000000000001000000000000001110100000000000010010000000000000001000000000000110000000000001101111111111111101111000000000001000100000000000010011111111111110111000000000001000100000000001011100000000000011110111111111111010011111111111001000000000000000001111111111110101111111111111100110000000000101001111111111111111100000000000110110000000000000110000000000001001100000000001011110000000000001011000000000000101100000000000100101111111111110101000000000001101000000000010100100000000001001010000000000001010100000000000011111111111111100011111111111111111111111111111110111111111111010111111111111111011011111111111101011111111111110000000000000001111000000000000000010000000000000000000000000000011000000000000010111111111111110100000000000001110000000000000000111111111111111100000000000010011100000000000001001111111111101100111111111111111011111111111011111111111111110010111111111101111011111111110010011111111111010010000000000000001100000000000010011111111111100100000000000000110111111111111111011111111111111001000000000000110111111111110111111111111111000001111111111111110000000000000001100000000000000000111111111111101100000000000001100000000000000100111111111101011111111111111011001111111111111110111111111110001100000000000001100000000000010010000000000000100000000000000011100000000000000000000000000000010000000000000011011111111111111100000000000000101111111111111110111111111111110010111111111110101100000000000001000000000000000001111111111111000011111111111100011111111111100011000000000000010111111111111111001111111111100100111111111111100000000000000111111111111111010001000000000010100000000000000100000000000000000101000000000000101011111111111011010000000000010001111111111110101111111111110111101111111111001111000000000000000011111111111110001111111111111010000000000001010111111111111101010000000000000000000000000000010111111111111010000000000000011011111111111110010111111111111001011111111110111000111111111111010111111111110111111111111111110111000000000000000000000000000000000000000000010001111111111111101011111111111110011111111111111110111111111111111011111111111110000000000000000010111111111101111011111111111100010000000000011001111111111111100011111111111100101111111111110011111111111111011111111111110101111111111111110000000000000000011011111111111001010000000000010001000000000001001111111111111010011111111111100100111111111111110111111111111010011111111111100101111111111111110011111111111010111111111111101010111111111111110000000000000101000000000000011100000000000001100000000000000000010000000000001100000000000000000111111111111101011111111111101010111111111110001100000000000000111111111111011111111111111111001000000000000011000000000000000000111111111111110111111111111111110000000000001000000000000000110111111111111111101111111111110111111111111111111111111111111011000000000000001101111111111111001011111111111011010000000000000000000000000011000000000000001101110000000000100001111111111111100100000000000010101111111111100001111111111110110000000000000000001111111111110110000000000000000011111111111101111111111111111001000000000000001111111111111101100000000000011011000000000000100011111111111110000000000000001111000000000010000000000000001101110000000000101101000000000001011000000000000011111111111111011110000000000001011011111111110110001111111111100111111111111111110100000000000011101111111111110110111111111110110111111111111010111111111111111101111111111111010100000000000000011111111111111001000000000000101111111111111110101111111111111101111111111111100100000000000000010000000000010111000000000000100100000000000110110000000000011110000000000100000000000000001011011111111111101111111111111111000000000000000001101111111111110111111111111111011100000000000000110000000000011010111111111111011000000000000011000000000000100011000000000010100100000000000011000000000000000111111111111111101000000000000001111111111111110010000000000011111100000000000100101111111111111101000000000000011000000000000101001111111111111100000000000000010011111111111110000000000000001001111111111111001100000000000010001111111111111110111111111111100000000000000100110000000000001010111111111111110011111111111101110000000000010011111111111111101111111111111110011111111111111010000000000000010100000000000000010000000000011001111111111110110011111111110111101111111111111110000000000000111011111111111111011111111111110000000000000001100111111111111111011111111111010000000000000100110000000000000101111111111111000101000000000000010111111111110101001111111111011011111111111011111011111111111001101111111111100110000000000010101000000000000101111111111111110011111111111111011011111111111111011111111111111101000000000000110100000000000010010000000000010011111111111111010100000000000010001111111111110111000000000001010100000000001101110000000000101100111111111111100011111111111111100000000000011100000000000000100011111111111000100000000000001010000000000010101100000000000001100000000000100010000000000000011100000000000000010000000000011110111111111110101011111111110110001111111111011001000000000001111111111111111111101111111111111010000000000001100111111111111111011111111111100001000000000010010100000000000101111111111110111100000000000000000100000000000110000000000000000001000000000000100100000000000000100000000000010000111111111101110100000000000010001111111111110000000000000000111000000000000001011111111111111001111111111110101011111111111100101111111111001011111111111111001100000000000111010000000000011001000000000001101111111111111011111111111111011010111111111111111000000000000101001111111111111100000000000010110011111111111101100000000000001100111111111111111000000000000000000000000000001011000000000000000011111111111011101111111111011100111111111111001011111111111110101111111111010001111111111101101111111111110111111111111111100111111111111110111100000000000000001111111111111101111111111111100100000000000011010000000000000111000000000000001100000000000001010000000000110110000000000000010000000000000101110000000000000001111111111111001111111111111101011111111111101100000000000000110100000000000101000000000000010001000000000001011111111111111101111111111111011011111111111110001111111111111111111111111111100101111111111111111100000000000000001111111111111011000000000010010111111111111111001111111111101101111111111110111000000000000011110000000000010110000000000010100000000000000000110000000000001010111111111111011111111111111010000000000000100001000000000001011111111111111111110000000000010100111111111101101011111111111001011111111111111111111111111111000000000000000011010000000000011110111111111111111100000000000001110000000000001000000000000000000111111111111011101111111111000001000000000010011100000000001011001111111111100110000000000010001011111111111110001111111111101011000000000001010111111111111110111111111111101100000000000010000000000000000010101111111111011111000000000001111011111111111110000000000000000101111111111110111111111111111011000000000000000100000000000000111100000000000110010000000000000110000000000000100100000000001100000000000000011100111111111111011011111111111110001111111111101100000000000011010111111111111110111111111111110110000000000010011000000000000011100000000000000101111111111111110100000000000001110000000000000111111111111111110000000000000010010000000000000011111111111111111011111111111001011111111111110101000000000001011000000000000010011111111111100101111111111111111011111111111111001111111111111100000000000000110100000000000001010000000000001000000000000000001100000000000000001111111111111010111111111111111000000000000000000000000000000101000000000001000011111111111110110000000000000000111111111110100011111111110100101111111111101111111111111101001111111111111001001111111111110000111111111111101011111111111001001111111111100110000000000000000100000000000000000000000000000000111111111111101100000000000001101111111111101011111111111110110111111111111110101111111111101011000000000000100111111111111101011111111111110111000000000001000100000000000001110000000000010000111111111111001100000000000110100000000000000011000000000000111000000000000001100000000000000001000000000000110011111111111010101111111111101110111111111110100011111111111100111111111111011110000000000000000000000000000010000000000000010100111111111111100111111111111011100000000000000001000000000001111100000000000011101111111111111010111111111111110111111111111110011111111111111100111111111111001011111111111101001111111111010001111111111111101100000000000011000000000000000001000000000001101100000000000101101111111111110010000000000000000100000000000001011111111111100111111111111100110111111111110101111111111111110110111111111111101000000000000010000000000000000111111111111111001000000000000011101111111111111100111111111111010111111111111101111111111111101110000000000000000100000000000000001111111111000011111111111110111111111111111100111111111111100011000000000000111100000000000100100000000000101010000000000001100100000000000010100000000000000000000000000001000000000000000100100000000000001010111111111111101011111111111101110000000000000110111111111111100011111111111011110000000000000000111111111111010011111111111000110000000000001010000000000000101000000000000100010000000000010010111111111111110000000000000111001111111111111111000000000000101000000000000110110000000000011010000000000000010100000000000011110000000000110001111111111111001011111111111100001111111111110000111111111110111100000000000000001111111111110010000000000000101000000000000110001111111111111010000000000000110000000000000000011111111111101111000000000000011100000000000000100000000000000001000000000000101100000000001001110000000000100110000000000010000000000000000101101111111111010100111111111110010111111111111100111111111111111001000000000000001111111111111100100000000000010101000000000000010111111111111111111111111111011100000000000000111111111111111111001111111111110101000000000010101100000000001100110000000000011100111111111100110011111111111011010000000000010100111111111110110011111111111011000000000000010000111111111110000111111111111100010000000000010000000000000011010100000000001100100000000000000100000000000010010100000000000011110000000000010010000000000000000111111111111110111111111111101101000000000000001111111111111011100000000000000000111111111111010011111111111101100000000000001011111111111111001011111111111100110000000000000000111111111111110100000000000001001111111111101010111111111111010100000000000000001111111111101100111111111110110011111111111110011111111111101011000000000010111100000000000101000000000000011101000000000000001111111111111011111111111111111011000000000000000011111111111001101111111111111110111111111111110000000000000100100000000000100000000000000000000000000000000010101111111111110110000000000001000111111111111110101111111111111000111111111111010100000000000010110000000000100110000000000010010011111111111110100000000000101000111111111111011111111111111101001111111111111111111111111110100100000000000010010000000000000001000000000000111111111111111110011111111111110010000000000000001111111111111111100000000000001011111111111110010111111111111100111111111111110100111111111111001100000000001001000000000000011011000000000001010000000000001011110000000000010110000000000000001011111111110111001111111111110111111111111111100111111111111000011111111111111001111111111111101000000000000000100000000000001101000000000000010000000000000000001111111111110101000000000000010011111111111101011111111111110010111111111111101100000000000000001111111111101110000000000000001011111111111101001111111111100110111111111110001111111111111111001111111111111110111111111111010011111111110101100000000000000000000000000001101000000000000111000000000000111010000000000000111100000000000010000000000000010111000000000000001000000000000110001111111111111100000000000000001111111111111100111111111111011110111111111110111111111111111001110000000000000010000000000001001000000000000010010000000000000001000000000000100111111111111011100000000000011101111111111111001111111111111001011111111111110100000000000000101111111111111101110000000000010010111111111111010100000000000100111111111111110100111111111111010011111111111010110000000000011001111111111111110000000000000001000000000000001000111111111111010000000000000100111111111110011111111111111111101011111111111100011111111111011111000000000000011000000000000001100000000000001111000000000001100100000000001000010000000000011110000000000000100111111111111110011111111111111110000000000000110100000000000010101111111111101001111111111101111011111111110011101111111111111101000000000000100011111111111110001111111111111111000000000000011100000000000001100000000000001100111111111111000000000000000010001111111111101000111111111111111011111111111110111111111111011101000000000001000100000000000100001111111111100011111111111110110111111111111101100000000000000010000000000001100100000000000011000000000000010001111111111111101000000000000011110000000000001101111111111110111011111111110000001111111111000101111111111110101011111111111001000000000000000010111111111111101100000000000001000000000000100010000000000000001000000000000000111111111111110011000000000000000011111111111001111111111111010111111111111110101111111111111101000000000000010110000000000010011000000000000001110000000000001011000000000001011000000000000100100000000000001100111111111111000011111111111000001111111111111100111111111111011111111111101010011111111111001101000000000001011111111111111101101111111111100100000000000001101100000000000001010000000000001111000000000000010000000000000011000000000000101001111111111111110111111111111011000000000000100001000000000010001111111111111111110000000000001100111111111111001000000000000100100000000000001111000000000000011111111111111110001111111111111011000000000000011000000000000000001111111111110011000000000001101011111111111110101111111110111111000000000000100100000000000000100000000000000110000000000001111000000000000110100000000000000111000000000000101100000000000010000000000000010011000000000001011100000000000010010000000000000000111111111111001100000000000001011111111111101111111111111101110111111111111001001111111111111000111111111111111000000000000101110000000000000101000000000000010000000000000101110000000000010101000000000000001011111111111110001111111111110101111111111111000111111111111100111111111111111010000000000000000100000000000101010000000000100010000000000001000011111111111110010000000000010000111111111111011111111111111101100000000000000100111111111111110111111111111101011111111111110010111111111110011111111111111110001111111111111101111111111111111111111111111010001111111111110010111111111111100011111111111100110000000000000001111111111110111111111111111011101111111111110010111111111111101011111111111100001111111111111101111111111111001111111111111101011111111111101100000000000000100000000000000000001111111111110101111111111111111100000000000000101111111111110001111111111110100100000000000001001111111111110101000000000000100011111111111110110000000000001001111111111111110111111111111111110000000000000010111111111111100100000000000100110000000000010100111111111101111011111111111101000000000000001010000000000000010011111111111111101111111111101011000000000000001000000000000011111111111111111110111111111110110111111111111110011111111111101111000000000000000111111111111010110000000000000010111111111110110000000000000110110000000000100110111111111111011111111111111100101111111111111010111111111110111011111111111011111111111111100111111111111111011100000000000000001111111111110111000000000000011011111111111101000000000000000000000000000001010100000000000000111111111111111000111111111111111011111111111101111111111111111001000000000000100000000000000010110000000000010101111111111111010100000000000000100000000000000111111111111110000011111111111011001111111111100110000000000000101100000000000111010000000000010101111111111111001000000000000101110000000000000111000000000000000011111111111100011111111111110111000000000000011111111111111111100000000000000111000000000000110100000000000111111111111111111111111111111111110011111111111011101111111111111111000000000000010000000000000001000000000000000010111111111111010011111111111101011111111111110010000000000000000111111111111010111111111111111101000000000000000111111111111000111111111111100101000000000000011011111111111111111111111111110011000000000000111111111111111111110000000000000001000000000000111100000000000010000000000000101001111111111111100100000000000101010000000000001101000000000000001100000000000000000000000000010011000000000001001000000000000001111111111111110010000000000000011011111111111100110000000000000010111111111111101111111111111110100000000000000010111111111111101011111111111100100000000000001110111111111110011111111111111111100000000000000010111111111111011111111111111101100000000000010100111111111111111000000000000000001111111111111100111111111111101011111111111111110000000000001110000000000000100111111111111111000000000000000101000000000001000000000000000010110000000000101101000000000000110100000000000101010000000000011111000000000001100000000000000011000000000000000110111111111111010100000000000011011111111111111110111111111111100100000000000000100000000000001000111111111111101000000000000010110000000000000100111111111111010111111111111101011111111111110100000000000000001111111111111101001111111111100001000000000001000000000000000000011111111111100000111111111110000100000000000001000000000000000000111111111111111000000000000101011111111111111100111111111111010011111111111101110000000000000000111111111111010011111111111100110000000000001011111111111111010111111111111111100000000000000000111111111111011100000000000011010000000000101010111111111110000111111111110010101111111111100001111111111111000111111111111011101111111111111011000000000000000100000000000011100000000000001100111111111111101111111111111100111111111111110010111111111111000100000000000010011111111111101000111111111110100000000000000100001111111111110100111111111111000111111111111001011111111111101110111111111110000111111111111011111111111111111010000000000011101100000000000100100000000000001101000000000000101011111111111110011111111111001111000000000000100011111111111111001111111111111010000000000010010100000000000100111111111111111101000000000001111011111111111111111111111111110011000000000000100011111111111100101111111111110110000000000000001000000000001001001111111111011000000000000000001000000000000001111111111111111100000000000000011011111111111011110000000000000100111111111110000011111111111001011111111111001100111111111110110111111111111110110000000000000011000000000001001000000000000000110000000000000000111111111110001011111111111100010000000000000001000000000000111000000000000100000000000000000101000000000000000100000000000101001111111111101000000000000000011000000000000000101111111111101001111111111111010100000000000000000000000000000000111111111111111100000000000000000000000000001000000000000010001100000000001001110000000000011100000000000000010011111111111011100000000000000101000000000000000011111111111110011111111111111000000000000000001000000000000001011111111111111110111111111111100011111111111011001111111111101111111111111110111011111111111100111111111111101010111111111110001011111111111100111111111111111100111111111110000111111111111000000000000000000101111111111111110111111111111000010000000000001110000000000001011100000000000000010000000000001010000000000001111100000000000001110000000000010011000000000000000011111111111111001111111111111011111111111111100111111111111100101111111111101010000000000001101000000000001011110000000000001011000000000000001111111111111101101111111111010101111111111111111100000000000010101111111111011100111111111110101011111111111111100000000000000110111111111111110100000000000000000000000000000000000000000000101000000000000011110000000000000100111111111110111111111111111101000000000000011110000000000000000000000000000011100000000000000000111111111111001000000000000001110000000000010101111111111111110011111111111011111111111111111101000000000000000111111111111010001111111111110001000000000000111000000000000011101111111111110111111111111111100011111111111010110000000000001000000000000000010111111111111101011111111111011111111111111101101111111111110010011111111111010000000000000001000100000000000111010000000000001101000000000000010000000000000011101111111111110011111111111111101000000000000001110000000000001010111111111110010011111111111000111111111111111000000000000000000000000000000000101111111111110101000000000010100100000000000100111111111111111001000000000000000100000000000010000000000000001111111111111111111100000000000011011111111111111011000000000000000100000000000010010000000000000001000000000000000100000000000000001111111111111001111111111111100100000000000001000000000000001110111111111111100011111111111010010000000000011101000000000000010100000000000010010000000000000000000000000100101100000000001001000000000000001000000000000000110000000000000001100000000000000101000000000000100100000000000111010000000000001110000000000000011011111111111111010000000000001111000000000010000100000000001000100000000000100010000000000011100100000000000110111111111111010011111111111110101111111111110101000000000000000010111111111111000100000000000111100000000000011100000000000000000000000000000110101111111111111010111111111111110000000000000000001111111111100111111111111111101011111111111111010000000000000011111111111111000000000000000100100000000000001011000000000000101000000000000011110000000000100101111111111111111011111111111101011111111111101010000000000010001100000000000000001111111111101100111111111111100111111111111001011111111111011010000000000000111000000000000100111111111111110011000000000001111100000000000000011111111111011110111111111110110011111111111010001111111111110101111111111111001000000000000100101111111111101001111111111111101100000000000001100000000000001001111111111111110100000000000000011111111111110000000000000001110011111111111111100000000000011110000000000000010000000000000001000000000000011011000000000000000011111111111100000000000000001010000000000001001011111111111101011111111111110101000000000000100100000000001000010000000000100010111111111111111000000000000100100000000000001100000000000000000011111111111111000000000000010000000000000010101000000000000000111111111111111000000000000000001100000000000011010000000000100101111111111110010011111111111010001111111111011010000000000000101000000000000011010000000000000011000000000000111111111111111101010000000000010000111111111111100000000000000001110000000000011000000000000010100011111111111101100000000000010111000000000000110111111111110111011111111111010100000000000000011011111111111110100000000000010000000000000000000000000000000000001111111111110001111111111111011011111111111010101111111111100011111111111111101011111111111001100000000000000110000000000001010100000000000000000000000000010001000000000000001011111111111011101111111111110011000000000000001000000000000001011111111111100011000000000001010000000000000001001111111111111011000000000010110000000000000001111111111111101110000000000000010111111111111111100000000000000011000000000000100011111111111110000000000000001011111111111111110111111111111100101111111111111011111111111101110011111111111111001111111111110001111111111110001111111111111101011111111111110101111111111110010011111111111110101111111111111100000000000001110100000000000001100000000000001001000000000001000100000000000010101111111111110001111111111111011011111111111101011111111111101000111111111101111111111111111101110000000000000110111111111101111111111111111000011111111111111000000000000000110111111111111011000000000000000101000000000001001000000000000000100000000000001010000000000000011000000000000101000000000000011100000000000000000011111111111100000000000000001010000000000000101111111111111101011111111111110100000000000000110011111111111001101111111111011101111111111110011111111111111100000000000000000000111111111110101000000000000011101111111111100111111111111111101011111111111101010000000000000000000000000000000100000000000000011111111111111011000000000000101011111111111101111111111111111011000000000000000011111111111010101111111111101110000000000000010000000000000010110000000000011000111111111111111000000000000010001111111111101010000000000000010111111111111111110000000000000110111111111111110111111111111111001111111111101101111111111111110111111111110101001111111111100111111111111101100011111111110011110000000000011000111111111110010011111111111100111111111111110101111111111111010111111111111000100000000000000011000000000000010000000000000101100000000000100010000000000011010000000000000010000000000000000010111111111111001111111111111010011111111111011101000000000000010000000000000001011111111111111001111111111111111100000000000101101111111111101011111111111111011100000000000000110000000000000001000000000100000000000000000011010000000000001010111111111110111011111111111100011111111111101000111111111111110000000000000011000000000000001011000000000010010111111111111100011111111111111010000000000001101100000000000100011111111111111111111111111110011111111111111101111111111111110000111111111111000100000000000000000000000000001000111111111111111111111111111011001111111111101100111111111111011111111111111011000000000000001001000000000000011000000000000000010000000000010010111111111111001111111111111100110000000000000000111111111111010011111111111100111111111111100111111111111101101111111111110111101111111111010010000000000001000100000000001000100000000000100010111111111111010000000000000010110000000000000101111111111110000111111111110110111111111110110110000000000000101100000000000011011111111111100101000000000001011100000000000010110000000000100010111111111111110000000000000110000000000000000111111111111111011111111111111101111111111111110001111111111110111111111111111100111111111111101000000000000000110011111111111101100000000000001100000000000000111011111111111010000000000000010100000000000000000011111111111110000000000000010000111111111011111111111111110011011111111111011011111111111111000111111111111110111111111111111101000000000010000011111111111011110000000000000000111111111111010011111111110111101111111111111001111111111110011111111111111010111111111111111010111111111110100000000000000000100000000000000000000000000000001011111111111111010000000000000001000000000000100000000000000101110000000000011101000000000000100000000000000011100000000000100010111111111110010011111111111110101111111111111111111111111111100100000000000011100000000000010011111111111111011000000000000100010000000000000010000000000000010000000000000111110000000000110000000000000000110100000000000011010000000000010100111111111111011011111111111011101111111111111000111111111111111111111111111111011111111111111010111111111111011100000000000000001111111111110101111111111111011100000000000000101111111111111000111111111110001111111111111010111111111111101010111111111101100011111111111111100000000000100001111111111111110000000000000100100000000000001101000000000000111100000000000000110000000000101010111111111101001011111111110111011111111111111101000000000001000100000000001000010000000000000110000000000000000011111111111101101111111111011010000000000001001000000000001011100000000000110001111111111110011100000000000001100000000000011000000000000001001000000000001000110000000000000000111111111101101011111111111100100000000000001000111111111100110011111111110110101111111111101101000000000001001000000000000001000000000000011111000000000000101111111111111111111111111111110110000000000000001000000000000000110000000000000110000000000001110100000000000011101111111111111101000000000000000000000000000011101111111111110001111111111110111111111111111100000000000000001111000000000000000011111111111101111111111111110100111111111110011111111111111000011111111111010010000000000000011100000000000110011111111111110100111111111111011111111111111000110000000000010001111111111110111111111111111110100000000000001011111111111101111111111111111110110000000000000110000000000000011000000000000110100000000000101000111111111110101011111111111100010000000000100101111111111101011111111111110101011111111111101100000000000001101000000000000010000000000000000100000000000001000100000000000001110000000000011000111111111111101000000000000001001111111111111010111111111111011000000000000100000000000000011101111111111111001000000000000100110000000000100011111111111101101111111111110101111111111111100110111111111111111111111111111011001111111111111110000000000001101100000000000011101111111111101001000000000000011100000000000110100000000000100101000000000010000000000000000110100000000000000000000000000001001100000000000011111111111111110001111111111111001011111111111110000000000000001110000000000000100011111111111111001111111111110101000000000000110100000000000011010000000000010111000000000001110000000000000010010000000000000101000000000000011011111111111011010000000000000110111111111111111111111111110101111111111111111010000000000000100011111111111110101111111111110101111111111101000011111111110011101111111111001000111111111111011111111111111000001111111111100110000000000001001111111111111110011111111111011001111111111110011000000000000001100000000000001000111111111111011100000000000001010000000000010000111111111110110000000000000000110000000000011011111111111111111011111111111010001111111111100001111111111111001100000000000001011111111111110010111111111111101111111111111100000000000000000101000000000001010000000000000110010000000000010010000000000000111000000000000001000000000000001110000000000000111011111111111111010000000000001000111111111111100100000000001001110000000000010101000000000000001100000000001000110000000000011101000000000000101100000000000011110000000000010001000000000000110011111111111010101111111111011000000000000001110111111111111111011111111111010011000000000000000000000000000000001111111111110000000000000010011000000000001000001111111111101101000000000010100000000000000001100000000000000110111111111110101111111111111110100000000000000110111111111111011111111111111001100000000000000001000000000000001100000000000000001111111111101000111111111111111011111111111010011111111111111100111111111110111100000000000000001111111111011100000000000001111100000000000010001111111111101011000000000001110011111111111000111111111111101100111111111111100000000000000001100000000000110101111111111111000100000000000100000000000000001111000000000000011011111111111001011111111111101110000000000000101100000000000011101111111111111111111111111111011111111111111011001111111111101000000000000000100011111111110111111111111111010111111111111111111111111111111110101111111111100110000000000001100000000000000011011111111111110001000000000000011100000000000000011111111111100100111111111110100011111111111101010000000000011000000000000000000000000000000000000000000000001111111111111101010000000000000001000000000000000100000000000000000111111111111011000000000000011101111111111111000011111111111100101111111111111101000000000000010011111111111111110000000000011101111111111110100100000000001001100000000000000101111111111101110011111111111111110000000000001001111111111110010111111111110101101111111111111110000000000000011000000000000000010000000000100011111111111111011000000000000000000000000000001110111111111111111100000000000011010000000000001110111111111111111111111111110100001111111111110100000000000000011011111111111110001111111111110001000000000000000011111111111110101111111111101001111111111111100100000000000000001111111111101010000000000010000100000000001100100000000000110110111111111110111111111111111010011111111111011110000000000001000011111111111111111111111111111110000000000000011100000000000001110000000000001011111111111111000111111111111111101111111111111111000000000000000000000000000111101111111111110100000000000000101111111111111100000000000000000100111111111111110111111111111010011111111111110111111111111110001011111111111110101111111111011101000000000001110011111111111101111111111111101110000000000001011011111111111111111111111111110100111111111111111111111111111110100000000000001100000000000000101100000000000100110000000000000001000000000000000000000000000000010000000000000101111111111111011011111111111100110000000000010011000000000000110111111111111101010000000000000111000000000000011111111111111101000000000000000000111111111110111000000000001100000000000000011010111111111111001011111111111101010000000000000100000000000000111111111111111011111111111111111011000000000000000011111111111001111111111111110100111111111111011011111111110111101111111111010101111111111111010100000000000000001111111111100110000000000000011100000000001001111111111111100110000000000000011000000000000001110000000000001000111111111111011111111111111111100000000000010100111111111111100100000000000100101111111111111100000000000000011000000000000000001111111111111010000000000000011011111111111111001111111111111000111111111101010011111111110010101111111111001101000000000000110000000000000110000000000000010011000000000001100000000000000100110000000000101000000000000000110000000000000000111111111111111010111111111111010100000000000001100000000000001001111111111111010011111111111110010000000000001010111111111110111111111111111010110000000000001111000000000000011011111111111101011111111111111000000000000000000100000000000010100000000000011010111111111111100111111111111001101111111111101100000000000000110000000000000100011111111111111101111111111111111000000000001011011111111111111111000000000001001000000000000001100000000000001111000000000000001100000000000011011111111111110101000000000001111000000000000000001111111111101010111111111110110100000000000001000000000000010111111111111111011100000000000000100000000000001101000000000001010111111111111110111111111111110111000000000010000000000000000000000000000000001001111111111110111011111111111101010000000000010101111111111111101111111111111110000000000000001000000000000000000000000000000000001111111111111111111111111111100111111111111010101111111111101111111111111111000111111111111011001111111111110101111111111110101011111111111100111111111111111001111111111110010111111111111111001111111111111001111111111110000111111111111101001111111111110001000000000000001111111111111101110000000000000111000000000000001011111111111110100000000000000001111111111111010011111111111101011111111111111101000000000001010011111111111110101111111111111010111111111111011100000000000001101111111111111111111111111111100111111111111110110000000000000110000000000000110000000000000101110000000000010110111111111111101000000000000010100000000000001111111111111111110011111111111010011111111111101011000000000000110000000000000010011111111111111111111111111110111111111111111010011111111111111000111111111110011000000000000110110000000000001001000000000000000100000000000011110000000000011010000000000000010000000000000001001111111111111011111111111110101011111111111111100000000000000011000000000001001111111111111101110000000000100011000000000000010000000000000100011111111111101110000000000001110000000000000110001111111111101101000000000000100100000000000000110000000000000011000000000000000011111111111111011111111111110110000000000000010100000000000010000000000000000110111111111111100011111111111001001111111111110010000000000001001011111111111011111111111111101101000000000001110011111111110111011111111111100001111111111111001111111111111000010000000000010101111111111101111011111111111011010000000000000000111111111101101011111111111110000000000000001110000000000001110100000000000000100000000000101000000000000000001011111111111010111111111111100110111111111101111111111111111010111111111111101000000000000000000000000000000101110000000000010100111111111110101000000000000000101111111111110101111111111111101011111111111111100000000000000100000000000010110100000000000101001111111111101110000000000010101000000000000001101111111111100100111111111111000000000000000101011111111111011010000000000000000011111111111011100000000000001000111111111111001000000000000110100000000000111011111111111111001100000000001011100000000000101010000000000000110011111111111100111111111111011110000000000001001011111111111101111111111111101000000000000001000000000000000010010000000000010000111111111111101011111111111111101111111111110011111111111111100111111111111101111111111111111111000000000000110100000000000100000000000000001101000000000000111011111111110110101111111111100111111111111110110111111111111011000000000000000110111111111101010011111111110101111111111111111001000000000001111000000000000101010000000000110100111111111110000111111111110110101111111111101011111111111111010011111111110110011111111111101001000000000000010100000000000101000000000001000000000000000000000000000000000001110000000000000000111111111110100100000000000000001111111111100110000000000001001011111111111101100000000000000010111111111110101111111111111000111111111111101000111111111110001111111111110101001111111111100100111111111110010111111111111101101111111111101000000000000000011011111111111011011111111111101101000000000000100100000000001000000000000000101111111111111100101011111111111101110000000000101011111111111101111100000000000000000000000000101010111111111111000100000000000101101111111111111011000000000000101011111111111111101111111111111000000000000001010100000000000000101111111111100110111111111111101111111111111110011111111111111100000000000010001100000000000000101111111111101110000000000010011011111111111111001111111111100001000000000000110000000000000000111111111111110011111111111100101111111111110110101111111111110001111111111110011011111111110011000000000000010000111111111111000000000000000010001111111111101111000000000001100000000000001001000000000000101100000000000001011100000000000101101111111111100001000000000000111100000000000000101111111111010011111111111111001111111111111101010000000000001001111111111111101011111111111110100000000000001110111111111111001111111111111111010000000000101011000000000010000111111111110110101111111111101001000000000000000100000000000001111111111111100011000000000000110111111111111011011111111111010101000000000001111000000000000000001111111111111111000000000000101011111111111011101111111111110011000000000000000100000000000000010000000000011100111111111101111000000000000000000000000000011110000000000000011000000000001010000000000000000100000000000000001000000000000110000000000000000000111111111100110111111111110110101111111111100110111111111110010000000000000001101111111111010011111111111101100000000000000011000000000000001011111111111111000000000000000000000000000000000110000000000000101011111111111111100000000000001011000000000000101100000000000110100000000000000100111111111111111111111111111010111111111111101100111111111111100011111111111100011111111111100010111111111101100111111111110111101111111111010000000000000001100111111111111100011111111111011011000000000001100011111111111100011111111111111011000000000001100111111111111111101111111111101000000000000001100100000000000001000000000000010111000000000001011111111111111101110000000000100011111111111111110000000000000101100000000000000000111111111111000000000000000010100000000000001000111111111110110100000000000000110000000000000111111111111111101100000000000001001111111111110110111111111101100011111111111101110000000000101011111111111101111111111111111110000000000000001101000000000000011100000000000000110000000000001101000000000001100011111111111111011111111110111010000000000001100011111111111011101111111111011000111111111110010011111111111000001111111111100011000000000000000111111111111111001111111111110111000000000000100011111111111100010000000000000100111111111110011111111111111110101111111111101001111111111111101111111111111111111111111111101011000000000000000011111111111110110000000000000000111111111111101111111111111110111111111111101101000000000000101100000000000110000000000000011110000000000000001100000000000010100000000000010101000000000011000000000000000011111111111111110010000000000010010000000000000001010000000000010110000000000000110000000000000001010000000000000111111111111111000000000000000111001111111111101100000000000000111111111111111101110000000000101001111111111111101000000000000000010000000000100111111111111111001011111111111101010000000000010010000000000000001000000000001001101111111111110111000000000000110000000000000100001111111111111011000000000000001111111111111100010000000000000000111111111110100111111111111100001111111111111100111111111111100000000000000011111111111111111111111111111111100011111111111110111111111111101011000000000001000011111111111111011111111111100100000000000000000111111111110100111111111111100110000000000001110111111111111010010000000000010110111111111110001011111111111100101111111111101101111111111110101011111111111100011111111111111000111111111110001111111111111100111111111111100011111111111101110011111111111110000000000000001100111111111110111000000000000010100000000000010010111111111111110000000000000111110000000000000100000000000001010100000000000001001111111111110010000000000000110100000000000010011111111111111010000000000000011011111111110010011111111111001001111111111110111011111111111101101111111111111011000000000000000011111111111101010000000000000110111111111110010100000000000000001111111111111101000000000000000100000000000011110000000000001101000000000000101000000000000000010000000000100001000000000000101011111111111101110000000000000001000000000010110000000000001100001111111111111100000000000000110011111111111001101111111111110101000000000000001011111111111101101111111111101110000000000000111100000000010001110000000000100001000000000001001100000000001110000000000000101011111111111111011100000000000010100000000000011111000000000000011111111111110110101111111111011000111111111111101111111111110101001111111111010100000000000000010011111111110101101111111111101011;
endcase
end
endmodule



module lut_weights_7(sbyte,addr);
input [3:0] addr;
output reg [124415:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0111: sbyte = 124416'b111111111111111100000000000011000000000000001011111111111111111111111111111111100000000000010111000000000000010111111111111100010000000000000111111111111111101100000000000100110000000000010001111111111111000100000000000000001111111111110000111111111101111011111111111101101111111111101011000000000001110000000000001011110000000000000010111111111110101011111111111100011111111111101101000000000000110111111111111010101111111111011101000000000010000000000000000001001111111111101011000000000000110011111111111111001111111111100101111111111101111111111111111101111111111111111100111111111111111011111111111110001111111111110001111111111111111000000000000100101111111111110101000000000001101100000000000000110000000000000000000000000011001000000000000101110000000000010011111111111111000100000000000000001111111111110010111111111110101111111111111000011111111111011000111111111111011011111111111101100000000000000101000000000001000111111111111100010000000000010100000000000000001011111111111011100000000000010100111111111110111000000000000001000000000000000000000000000000100011111111111011010000000000000000111111111111110111111111111111110000000000010000111111111111100100000000000011101111111111111110000000000000001000000000000001000000000000011110111111111110010100000000000110101111111111111111111111111111011011111111111100111111111111111101000000000000101011111111111101010000000000000100111111111111000011111111111101101111111111100100111111111111100100000000001001111111111111110010111111111110111011111111111110000000000000000110111111111111000100000000000000011111111111111100000000000001011000000000000000110000000000000010111111111111111100000000000000000000000000000111000000000000111100000000000010110000000000000001000000000011000100000000000010000000000000000000000000000010101111111111111101110000000000000000000000000000001100000000000011001111111111100100000000000010010100000000001010110000000000011000000000000000100000000000000000011111111111111101000000000000111100000000000001111111111111001010111111111111011111111111111111011111111111110100111111111111110111111111111111101111111111111011000000000000000111111111111001000000000000000011000000000001010000000000000001000000000000001011000000000000111100000000000000100000000000001110111111111111000111111111111111111111111111111101111111111111110011111111111111011111111111110111111111111111011011111111111111001111111111111101111111111111111100000000000010100000000000010111111111111110011100000000000001111111111111110011111111111111100011111111111001110000000000001001111111111111000000000000000000111111111111110111111111111101000111111111111100010000000000011101000000000000000100000000000000011111111111110000000000000000010000000000000000001111111111111101111111111110110011111111111101000000000000000000111111111111110111111111111000100000000000010100111111111110100111111111111100100000000000000010000000000000101000000000000001100000000000010001111111111110101111111111111111110000000000001000000000000001001011111111111110011111111111111101000000000000011100000000000100100000000000001110000000000000011000000000000001000000000000011001111111111111111100000000001000010000000000000001000000000000000011111111111101000000000000001011000000000001001011111111111110101111111111111010000000000000001111111111111000101111111111101001000000000001111011111111111000001111111111110011000000000010010000000000000001011111111111100110000000000001001000000000000100110000000000100011111111111111001000000000000011010000000000000001111111111111000111111111111101011111111111111010000000000000000111111111111110011111111111110110111111111111101011111111111110010000000000100001111111111111110000000000000100001111111111110100000000000000111100000000001000001111111111110000000000000000000000000000000110010000000000011101000000000001001011111111111101001111111111101110000000000000001100000000000010110000000000000111000000000001010100000000000111011111111111100110111111111111110000000000000000101111111111111111111111111111110100000000000001001111111111111101111111111111010000000000000011100000000000000000000000000000101000000000000001000000000000000011000000000000011011111111111110011111111111110110000000000000100100000000000010011111111111111001111111111111010111111111111010011111111111111111000000000000000000000000000000011111111111101000000000000001011000000000000000000000000000010000111111111110101111111111111101011111111111101111111111111110001111111111111110011111111111111110111111111111001100000000000100110000000000001001111111111111100011111111111101001111111111111101111111111111100011111111111111010000000000001100111111111111001011111111111111100000000000010010000000000000100111111111111010101111111111111111000000000000001000000000000000110000000000011100000000000000011000000000000000001111111111100101111111111110110000000000000000100000000000010011000000000000000100000000000010100000000000001001111111111111100111111111111110001111111111110001000000000000001000000000000000001111111111101000000000000000010111111111111111011111111111100011000000000001010100000000000101111111111111101001111111111111011100000000000100100000000000001000111111111111010111111111111110111111111111110011111111111111110000000000000000000000000000000000000000000000001000000000000011000000000000010101000000000000101000000000000010101111111111110111111111111111101011111111111111100000000000011010000000000001000000000000000001110000000000000111111111111110100100000000000001100000000000001111111111111111110011111111111101111111111111110101111111111111010111111111111111111111111111110001111111111111011000000000000000101111111111101010000000000000001000000000000000000000000000000011000000000001001000000000000110010000000000010000000000000001111100000000000000001111111111011100000000000001001011111111111101010000000000001001111111111111111111111111111001010000000000010110000000000000010011111111111100100000000000000000111111111110111111111111111111100000000000000110111111111111011011111111111111001111111111110000000000000000010111111111111010010000000000000011111111111111000011111111111000100000000000001001000000000000101000000000000001100000000000001101111111111111000011111111111010000000000000001010111111111111110011111111111110001111111111110001111111111111001111111111111010010000000000010110111111111110111100000000000000011111111111110100111111111111111000000000000010010000000000000101111111111110110011111111111111000000000000001100111111111110101000000000000111110000000000000011111111111110100100000000000101011111111111110100111111111111000111111111111110111111111111110100111111111111100011111111111111001111111111111011111111111111100000000000000001101111111111001101000000000000000000000000000010010000000000001110000000000010011011111111111111001111111111010011000000000000011111111111111110111111111111110010000000000001010011111111111010101111111111100010111111111110110011111111111111110000000000001001000000000000000000000000000000001111111111101110111111111111111011111111111011100000000000001111000000000000010100000000000010101111111111101101000000000000010000000000001011011111111111111101111111111111100011111111111101110000000000001101111111111111000011111111111010001111111111011010000000000011001000000000000111000000000000111101000000000010111100000000001111001111111111110100000000000000100011111111111001001111111111100110000000000000111000000000000111000000000000001001111111111111001000000000000000111111111111110001111111111101100111111111111010000000000000000000000000000000000000000000001000111111111111011100111111111111101100000000000101111111111111011011111111111111010011111111111010011111111111110000000000000000001000000000000010010000000001100011000000000000110000000000000010101111111111011001111111111101111111111111110101011111111111011000111111111111011111111111110111011111111110101011111111111111101011111111110111011111111111101101111111111110000011111111110111110000000000101010111111111111110111111111111110111111111111111010111111111110111011111111110111111111111111111000000000000000101111111111111110100000000000001110000000000000000000000000000101000000000000000001000000000000001100000000000001010000000000010111111111111111001011111111111000010000000000000000000000000000011011111111111101000000000000000001111111111111000011111111111001100000000000000001111111111111111000000000000101011111111111101000000000000001011011111111111011001111111111101001000000000000011111111111111111001111111111101111000000000000000011111111111100011111111111110011000000000010101000000000000101111111111111101010111111111111001011111111111001111111111111111011111111111111010011111111111010101111111111101011000000000010010111111111111100111111111111010101111111111111101100000000000101000000000000100100000000000001000000000000001000001111111111110111000000000010010000000000000110000000000001000001111111111110100111111111111111100000000000000101111111111110100111111111111010111111111111101000111111111101110011111111110101011111111111001010000000000000110000000000000110100000000000010010000000000000010111111111111001001111111111110110000000000011101100000000001001110000000000010001000000000000111111111111111110100000000000100110000000000001110011111111111111111111111111100100000000000000011100000000000000001111111111101001000000000001000000000000000001111111111111111000000000000001010111111111111100000000000000010110000000000000011111111111111001101111111111101000000000000000100000000000000001100000000000000000000000000000011111111111111011001111111111101001111111111101111111111111110011001111111111110101000000000000001100000000000010101111111111111001000000000001010100000000000100100000000000000111111111111110110011111111101100111111111111101100111111111100101011111111110001000000000000001010111111111101110011111111110101101111111111111001000000000001011000000000000111110000000000000010000000000001000111111111101111111111111111110111000000000000110100000000000011101111111111101110000000000001110100000000000010101111111111100100000000000001000011111111110100011111111111101111111111111110011111111111111010001111111111100111000000000011001000000000000000011111111111111111111111111111100000000000001001101111111111111110000000000001100000000000000110111111111111101111000000000000111100000000000010101111111111111001000000000000001011111111111011011111111111101111111111111110100011111111110111010000000000000111111111111111110100000000000110111111111111111101111111111111110011111111111110100000000000010110000000000000101011111111111011110000000000000001000000000000000111111111111010110000000000000000000000000001111111111111111100111111111111110000111111111110110111111111111010011111111111101010000000000010010100000000000000101111111111111010111111111110010100000000000000111111111111110101111111111111000100000000000100111111111111111101000000000000110011111111111110011111111111100111000000000000011111111111111111110000000000000101111111111110100011111111111110110000000000010000000000000011001011111111111110111111111111111101000000000001010000000000000001111111111111111001111111111111110111111111111100000000000000010110000000000000100111111111111110110000000000010000111111111111011111111111111011100000000000000000111111111110000111111111111001001111111111100101000000000001011100000000001000110000000000010000000000000001101000000000000011000000000000001111000000000000000000000000000010110000000000000101000000000000010011111111111111001111111111111110111111111111111100000000000001100000000000001001111111111111001000000000000000100000000000000011111111111111010111111111111100100000000000000100000000000000100000000000000011100000000000001010111111111111100011111111111010110000000000000001000000000000101000000000000001110000000000011011000000000001011111111111111110100000000000001100000000000000000011111111111111011111111111111011111111111111001011111111111001000000000000001111111111111111110000000000000110001111111111111010000000000000101000000000000101000000000000001011000000000000011100000000000000110000000000011100111111111111000100000000000010100000000000001111000000000000011011111111111011100000000000000100000000000010100100000000000010011111111111010101111111111111010111111111111111101111111111100000111111111111101011111111111010110000000000001110000000000010110100000000001010011111111111111001000000000000100111111111110111111111111111101000111111111111101011111111111101101111111111100111000000000000011000000000000110100000000000010101000000000000110011111111111111001111111111111101000000000000001100000000000101000000000000000000000000000000100011111111111100101111111111010110000000000000010011111111111001111111111111111100111111111110111011111111111100010000000000001101111111111111100011111111111111101111111111111111000000000000101100000000000001010000000000000000000000000000010111111111111111011111111111111101111111111111101000000000000011010000000000001110000000000000110100000000000111110000000000000111111111111101111111111111110111001111111111101010111111111110011100000000000000001111111111110011000000000000110000000000000101011111111111110011000000000001111000000000000011010000000000000001000000000000110100000000000100000000000000001010000000000000111011111111111111001111111111110000111111111111100111111111111010101111111111111110000000000000111011111111111101110000000000001111111111111111111000000000000010000000000000011000000000000000100000000000000101111111111111101010000000000000011000000000000011100000000000000100111111111111011100000000000111011111111111111001000000000000100111111111111100011111111111101100000000000000010000000000000000011111111111110110000000000000110100000000000010011111111111110000111111111111010011111111111110011111111111110101111111111111111111111111111100101111111111110000111111111111001000000000000011110000000000011010000000000000010000000000000011001111111111111101111111111111011011111111111000111111111111110010111111111111111111111111111110111111111111111100000000000000011011111111111101110000000000010010000000000000101000000000000001001111111111011111111111111110010111111111111010101111111111111011111111111101001111111111110111111111111111110101000000000001111011111111111110000000000000011010000000000001101111111111111110100000000000001011111111111111000011111111111110001111111111100001000000000000100000000000000101000000000000000111000000000001001111111111111010111111111111110001111111111110010111111111110101111111111111100101000000000010100000000000000011000000000000001110000000000000011111111111111101111111111111111001111111111111110011111111111001011111111111011101000000000001101100000000000001100000000000011110000000000000010100000000000000001111111111111100111111111110010011111111111110010000000000000000111111111111100111111111111111001111111111110111000000000001000000000000000100010000000000010000000000000001010000000000010001001111111111111110111111111110110011111111111101111111111111110110000000000000011000000000000100010000000000000001000000000001101011111111111111000000000000000101000000000001111100000000000110011111111111101001000000000001110100000000000010101111111111111001111111111110101111111111110100011111111111010111000000000001100011111111111111001111111111011110111111111110101011111111111110100000000000001001000000000000000000000000000010000000000000010111111111111111010111111111111001101111111111111101111111111111111111111111111110110000000000000010000000000000100100000000000011000000000000000100000000000001111011111111111010001111111111011010111111111111100111111111111001011111111111111011000000000000000011111111111110101111111111101100000000000011011111111111111111111111111111111011000000000001010111111111111100010000000000000000000000000001100000000000000000100000000000000101000000000101000011111111111101111111111111100001111111111110100100000000000000101111111111101110111111111111001100000000000101001111111111101110000000000000101111111111111100011111111111111111000000000000101000000000000101000000000000010110000000000001001011111111111011111111111111100100000000000001100111111111111011100000000000100000000000000000100100000000000001010000000000001001000000000000000011111111111111001111111111101101000000000001000111111111111111110000000000001100000000000000100000000000000010010000000000000101000000000000100100000000000101011111111111110101111111111101110111111111111010111111111111100011000000000000111000000000000001001111111111111111111111111111101100000000000000011111111111111001111111111111011111111111111011011111111111110110000000000000001111111111111100101111111111111110000000000001110000000000000100111111111111101110000000000000101011111111111100111111111111101011111111111111000011111111110101110000000000001010111111111110011111111111111010011111111111111000111111111110000100000000000001010000000000000010000000000000000100000000000001111111111111101111000000000010100000000000000100111111111111111010000000000001100000000000000100101111111111110000000000000000001111111111111100110000000000000001111111111111010011111111111110100000000000001101000000000001110111111111111101000000000000011010111111111111111000000000001000010000000000000000000000000000110000000000000010010000000000000100000000000000100011111111111111011111111111110011000000000001100100000000000000001111111111110101000000000000111000000000000110110000000000000000000000000000101000000000001001001111111111111100111111111110101011111111111101100000000000000100111111111110100100000000000000010000000000010011000000000010110011111111111010111111111111100001000000000010100100000000000001100000000000010000111111111111100011111111111011110000000000000000111111111111111111111111110011111111111111101001000000000000100011111111111111111111111111111101000000000000100000000000001010111111111111111010000000000000010100000000000110000000000000100000111111111111100111111111111111100000000000010011111111111101111011111111111001101111111111110010000000000000000000000000000100000000000000110011111111111111111111111111111011110000000000000101000000000000010000000000000101000000000000001010000000000000001011111111111011101111111111111110111111111111011000000000000101000000000000110010111111111101110011111111111000000000000000001111111111111110011011111111111011111111111111111001111111111111111011111111111111011111111111111101000000000001011000000000000000000000000000000000111111111111010111111111111110110000000000000011111111111110110000000000000110010000000000001001111111111111001000000000000100100000000000000010000000000000001111111111111111110000000000011010000000000001100111111111111110110000000000001100111111111110111000000000000000111111111111001010000000000000111000000000000011111111111111100001000000000001110000000000000011010000000000001010111111111110001011111111111001110000000000011000000000000000001000000000000001010000000000000101111111111110101100000000000101101111111111111111111111111110001011111111111110011111111111011111111111111111100111111111111010111111111111101011111111111111001011111111111010101111111111101101000000000000001100000000000111100000000000010101111111111110110100000000000101101111111111111110111111111111100111111111111011001111111111111101000000000001010111111111111111110000000000000001111111111111011011111111111010011111111111101000000000000001110000000000000100011111111111101110000000000010010100000000000011100000000000000010000000000000110111111111111111100000000000000000000000000000010100000000000000111111111111111110111111111110000000000000000011110000000000010000111111111110111011111111111111011111111111110010000000000000000011111111111100110000000000001101000000000001010011111111111101100000000000011100000000000000010111111111111110111111111111110100111111111111101000000000000110000000000000001110000000000000010100000000000000100000000000100101111111111111000111111111111110101111111111111101000000000001010100000000000001001111111111110000000000000000000011111111111010011111111111101001000000000001010011111111111101111111111111110010000000000000010111111111111111101111111111111110000000000000110000000000000010000000000000001000111111111111110100000000000101100000000000011100111111111111111011111111111111110000000000001000000000000000010111111111111100001111111111101001111111111101100011111111111011110000000000101010000000000000000011111111111010101111111111111111111111111111111100000000000011111111111111110100111111111111011011111111111101101111111111111100111111111111001000000000000001101111111111111111000000000000101000000000000101000000000000000100111111111111001111111111111100000000000000001011111111111111111111111111111111110000000000000010000000000000000011111111111000100000000000100101000000000001000111111111111111000000000000000001000000000000000100000000000011000000000000001100111111111110001100000000000001010000000000010011000000000000010100000000000000001111111111101010000000000000100111111111111110011111111111111010000000000000010100000000000000110000000000000110111111111110101100000000000000001111111111001110000000000000000011111111111011000000000000011110000000000000110000000000000110100000000000100000111111111111111011111111111111011111111111111110111111111111100100000000000000100000000000001110000000000000011000000000000100010000000000001100000000000000111000000000000011100000000000010011111111111111101111111111111010010000000000001100000000000001001100000000000001100000000000000001111111111111100100000000001000100000000000001010111111111111111111111111111101001111111111011101000000000001100000000000000001000000000000001010111111111111111100000000000001000000000000000101111111111111000111111111111011111111111111100111000000000001011000000000000101110000000000000111111111111111110000000000000010111111111111111111000000000000000111111111111111111111111111011010111111111111010111111111111001011111111111101001111111111111011000000000000000110000000000001111000000000000010100000000000110000000000000000000000000000000010011111111111110101111111111111011000000000000001000000000000000001111111111101000000000000000011011111111111111001111111111111011000000000010001100000000000100110000000000100010000000000000011011111111111001011111111111110111000000000000000111111111111101000000000000010110000000000000001111111111111110111111111111010111111111111111010111111111110100111111111111101100000000000000011100000000000000100000000000011100111111111111101000000000000001000000000000001111000000000001100011111111111100001111111111111011000000000001101000000000000000001111111111111100000000000010100111111111111100000000000000001110111111111110101111111111111011001111111111100100111111111110101100000000000100010000000000101110000000000000000100000000000100011111111111110110111111111110110111111111110110010000000000001001111111111111000000000000000011000000000000001110000000000000111000000000000001011111111111110000111111111110011100000000000010011111111111101100111111111110110000000000000000110000000000011010000000000001011100000000000010010000000000000000111111111111011011111111111110011111111111101100111111111110110000000000000001100000000000101010111111111111100111111111111110001111111111101001000000000000011000000000000000110000000000001010000000000000000000000000000010011111111111110110111111111111110100000000000001101111111111111111000000000000101100000000000000000000000000001111000000000000100000000000000001111111111111111101000000000000001111111111111100001111111111110111111111111110100000000000001000001111111111111110000000000000011111111111111100100000000000001101000000000000010000000000000000000000000000001110000000000001101011111111111101101111111111111001111111111111111100000000000000000000000000000000000000000001000011111111111111010000000000010001111111111111001011111111111101001111111111101101111111111111011011111111111111000000000000010001111111111111101000000000000011010000000000010101000000000000011000000000000000001111111111111100111111111111100100000000000000001111111111111100111111111110111100000000000010010000000000000011111111111111001011111111111101111111111111111100111111111110101100000000000011010000000000010100000000000000000100000000000001101111111111111111000000000000110100000000000110000000000000011100111111111111011100000000000001000000000000010100000000000000010100000000000101001111111111111111000000000000110011111111111111111111111111100110000000000000001111111111111110111111111111110010000000000000001100000000000100001111111111111010000000000001110000000000000101100000000000001101000000000000100100000000000100001111111111010000000000000001001000000000000001001111111111100011000000000000011100000000001000101111111111111110111111111111001011111111111011000000000000000001000000000001101011111111111110001111111111111101000000000010111100000000001001001111111111100001111111111110000011111111111111011111111111001111000000000000011000000000000101010000000000010000000000000000000011111111111000010000000000011100111111111111101000000000000011011111111111110011000000000000001111111111111110001111111111110001000000000001100100000000000110101111111111001011111111111111100100000000000011111111111111101011000000000001110111111111111110100000000000010110111111111110001111111111111101100000000000000111111111111111101011111111111011110000000000001110111111111110100011111111111111000000000000010111111111111111011100000000000011100000000000000110000000000001010111111111111010001111111111111100111111111111000100000000000001001111111111111100111111111110111100000000000000100000000000010100111111111101010011111111111111111111111111111101111111111111000100000000000011000000000000011111111111111101111111111111111010001111111111111010111111111111100000000000000110010000000000010010000000000001100100000000000000011111111111100101000000000001100100000000001101001111111111110000111111111111101011111111110111011111111111101010000000000010000011111111111101110000000000000100111111111111110100000000000110100000000000100100111111111111001000000000000011110000000000000000111111111111010000000000000000110000000000000001111111111110001111111111111010100000000000101100000000000000001100000000000011110000000000010111000000000010000000000000000100001111111111111101000000000000101000000000000101000000000000001110111111111110000111111111111111000000000000010010000000000000011111111111111101001111111111110110111111111101000111111111110110100000000000010001111111111110100111111111111001111111111111111000000000000000001011111111111100000000000000001101111111111100110111111111111011000000000000110000000000000001001000000000000100011111111111101011111111111111010111111111110110100000000000010111000000000000010111111111111010010000000000001101111111111111001111111111111101000000000000001101000000000000110000000000000000000000000000000100111111111111101111111111111110100000000000001000000000000000010011111111111010011111111111101011111111111110111100000000000111010000000000010011000000000001001100000000000010110000000000001101000000000001010011111111111011100000000000000111111111111101110111111111111001111111111111110001000000000000110100000000000101111111111111110001111111111101100100000000000100010000000000010110111111111111000100000000001001000000000000011100111111111111111111111111111110000000000000000101111111111110110100000000000001100000000000001001111111111111000011111111111110001111111111000100000000000000011000000000000000010000000000011001111111111110111000000000000111010000000000000010111111111110100000000000000010000000000000100000111111111101110111111111110111011111111111110000000000000001101111111111111001001111111111011110000000000001000100000000000101011111111111001010111111111101101111111111111000100000000000011000111111111110111011111111111101101111111111111001111111111111010000000000000001000000000000001100111111111111110100000000000000011111111111101001000000000000100100000000000001001111111111111001111111111110100000000000000100101111111111110011000000000001001011111111111110010000000000000101000000000000100011111111111110100000000000000000000000000001010000000000000011001111111111101011000000000010010100000000000100100000000000000100000000000000110000000000000001011111111111111100111111111101111011111111111111000000000000000001000000000001001111111111111100000000000000001110000000000001010100000000000111000000000000010001000000000000000100000000000001010000000000010000000000000000011100000000000000000000000000000000000000000001110100000000000001110000000000100011111111111111000011111111111101000000000000001010000000000000010111111111111100101111111111101110111111111111011111111111111100101111111111111111000000000001001000000000000000000000000000000110111111111111000111111111111101000000000000000110000000000000100011111111111110101111111111011101111111111110100111111111111111101111111111100001000000000000011111111111111111110000000000100011111111111111110011111111111010010000000000000010111111111111010011111111111111100000000000010001000000000000111011111111111110000000000000011101000000000000101011111111111110010000000000000111111111111111110011111111111011010000000000001011000000000000011000000000000110101111111111100111111111111111101111111111111011011111111111100110111111111111111100000000000001001111111111111000111111111110001000000000000000001111111111110011000000000000101011111111111101111111111111101001111111111111100111111111111100010000000000000000000000000000111011111111111110000000000000010010000000000001111100000000000111011111111111111100111111111111001011111111111001100000000000001001000000000010000000000000000111011111111111101100111111111111110000000000000110101111111111100111111111111111100100000000000000001111111111111000111111111111000000000000001001001111111111110001111111111111100000000000000001010000000000000011000000000000100011111111111000010000000000100001111111111111110100000000000111111111111111111010000000000000011111111111111110100000000000001110000000000001001000000000000001001111111111101001000000000000111111111111111010111111111111010011000000000000010111111111110111101111111111110000000000000001111000000000000001110000000000010011111111111111101011111111111010110000000000011010111111111111100100000000000011010000000000001001111111111111110000000000000010110000000000011100000000000000110011111111111101010000000000000011111111111111010111111111111111111111111111110010000000000000100000000000000011110000000000101001000000000000110111111111111001110000000000010111000000000000011111111111111111101111111111110111111111111111010011111111111110000000000000000000000000000001101111111111111111101111111111101110000000000000000011111111111111101111111111110111000000000000000011111111111100001111111111110001111111111110011111111111111011000000000000101010111111111111101100000000000001101111111111110010111111111110111111111111111111100000000000011101000000000000010000000000000111011111111111111000111111111111001100000000000011011111111111110110111111111101111100000000000000011111111111110101111111111111101100000000000010101111111111101000000000000001001111111111111111111111111111011010000000000010101100000000000010101111111111111001000000000000000011111111111100110000000000100011000000000000011100000000000000000000000000101001111111111111010011111111111110010000000000000001000000000001011000000000000100000000000000000100111111111101100011111111111111100000000000001101111111111111110100000000000101000000000000001101000000000001001000000000000000001111111111111011000000000100001000000000000101110000000000001010000000000000010011111111111011010000000000000000111111111111010000000000000100101111111111101000000000000000100000000000000100001111111111111110111111111111101100000000000000110000000000001100000000000001111111111111111110111111111111101000000000000010011000000000000111010000000000001100111111111111100111111111111011101111111111100000000000000000111000000000000101110000000000100101000000000000000011111111111111000000000000000011111111111100110011111111111010001111111111101000000000000001000011111111111010101111111111100111111111111111001111111111111111110000000000010010000000000000111100000000000000110000000000100110000000000001010000000000000100110000000000100001111111111110101000000000000101011111111111110111000000000011011100000000001001000000000000011011111111111111011111111111111100011111111111110100111111111111000111111111111101100000000000010011111111111111011111111111111001001111111111111001000000000000101111111111111101000000000000000111000000000001100100000000000000011111111111101110111111111101011111111111111100001111111111110110111111111111101100000000000000101111111111101011000000000000101100000000000010100000000000001011111111111111111100000000000000010000000000100101111111111110000111111111110110111111111111001111000000000010101000000000000011110000000000011000000000000001101100000000000010100000000000010111111111111111011100000000000100010000000000000001000000000000000000000000000101101111111111111000111111111110000011111111111111011111111111111001000000000000110011111111111010001111111111001100000000000000000011111111111100101111111111100101000000000001001100000000000010000000000000001010000000000001101011111111111111111111111111011010111111111111000100000000000001100000000000100110000000000000001011111111111111100000000000100100000000000000101100000000000100010000000000011001000000000000001011111111111000101111111111101100111111111111110111111111111010101111111111010010111111111111001011111111111101001111111111001110111111111101110100000000000000111111111111100111000000000001001000000000000001010000000000101000000000000000111000000000000101100000000000001010000000000000000011111111111101101111111111111010000000000001001100000000000000011111111111110001000000000000000011111111101110111111111111110111000000000001011011111111111011111111111111110101000000000011011100000000000110110000000000000110000000000001000011111111110101101111111111011101111111111111100011111111111111100000000000001001111111111111001111111111111111101111111111111110000000000001011000000000000011000000000000011100000000000001110000000000000100010000000000000011111111111110010111111111111111100000000000000101000000000001011000000000000110110000000000100111111111111110110111111111110101111111111111001110111111111111010100000000000110001111111111111101000000000000000100000000000101101111111111110100000000000001010100000000000111011111111111110011111111111101101000000000000010011111111111111101000000000000011000000000000000001111111111111000111111111101011111111111111010111111111111110101000000000001110100000000000100000000000000011111111111111101000111111111111000011111111111001010000000000000001100000000000010101111111111111110111111111111011011111111111101000000000000010101000000000001000000000000000010000000000000000001111111111101111100000000000001101111111111101101111111111111110011111111111101100000000000001000000000000000000011111111111011101111111111111100000000000001101011111111111101110000000000100000111111111111010111111111111010000000000000000000111111111111110011111111111110101111111111111101000000000000010111111111111110010000000000010101000000000000101100000000000000001111111111111001000000000001001011111111111111110000000000000101111111111110100100000000000110100000000000001100111111111111010011111111111010000000000000010000000000000000000000000000000000011111111111011011000000000000010011111111111111001111111111101011000000000000000111111111111100111111111111101111111111111110010111111111111111011111111111010001000000000000011100000000000110011111111111101000111111111110111000000000000100010000000000000110000000000000010000000000000011110000000000001110111111111111001011111111111011110000000000000111111111111111111011111111111100100000000000110110111111111111101111111111111101111111111111111100111111111111111000000000000001001111111111111010111111111110000100000000000000001111111111110101111111111110111011111111111110011111111111100111111111111110110011111111111110000000000000000000111111111111100100000000001011000000000000100011000000000000010000000000000001000000000000010011000000000010001100000000000011111111111111011110111111111110111111111111111101011111111111101101111111111110010111111111111101010000000000001011111111111111001100000000000010110000000000011010111111111111010011111111110111111111111111101001000000000000000011111111111101111111111111011110111111111110011011111111111100010000000000001010000000000011001100000000001010000000000000011101111111111110010011111111111011010000000000000010111111111110101000000000000001011111111111111100000000000001010111111111111101111111111111101100111111111111010111111111111100101111111111110111000000000000110111111111111101111111111111111000000000000010111100000000001011110000000000000001111111111111100000000000000000000000000000000011000000000000010100000000000100001111111111110000111111111110111111111111111010000000000000000110111111111100111111111111110110111111111111110101111111111110111111111111111110011111111111100101111111111101111111111111111101101111111111110101111111111111100011111111111110101111111111110101000000000001000000000000000001110000000000000011000000000000101111111111111110110000000000100011111111111111110011111111111100010000000000000111000000000010000111111111111001010000000000000001000000000010011011111111111110101111111111110101111111111111100111111111111101110000000000000011000000000000111111111111111111101111111111111101111111111111011111111111111111000000000000001100111111111111110011111111110100010000000000000111000000000000000100000000000000000000000000000000111111111111101111111111111000001111111111111110111111111111100100000000000001011111111111011110111111111111001100000000000000001111111111110101111111111110011100000000000101001111111111110110000000000000000111111111111111011111111111101001111111111111011111111111111011010000000000010111000000000001101100000000000010001111111111110000000000000000001111111111111011011111111111111100000000000000000100000000000110011111111111110111111111111110100111111111111111100000000000001100111111111111101000000000000001001111111111100011111111111110010011111111111101010000000000000000111111111111111000000000001011000000000000010011000000000000110111111111111100111111111111101111000000000000000011111111111100100000000000000101111111111111101100000000000000000000000000001000000000000001010000000000000001100000000000010101111111111111010100000000000001001111111111101000111111111110110000000000000000110000000000000000000000000000000011111111111001010000000000010001000000000000010000000000000010010000000000000110111111111110111000000000000100110000000000001010111111111111111111111111111100011111111111111110000000000000010000000000000001100000000000000000000000000000100000000000000000101111111111100011000000000001001111111111111110110000000000110110000000000000100100000000000011001111111111100001111111111111000100000000000100001111111111111111000000000000011011111111111110010000000000000010000000000000111100000000000011100000000000001100111111111111101000000000000000110000000000001011000000000000010011111111111110011111111111100011000000000000100011111111111100100000000000011010000000000001001000000000000101010000000000001011000000000000110000000000000010010000000000000001000000000000000111111111111111111111111111111011111111111111101000000000000000000000000000000001111111111111011000000000000001101111111111111010000000000000010000000000000001101111111111101000111111111111010100000000000000111111111111110001111111111111110111111111111101100000000000000111111111111110111000000000000000001111111111101000111111111111111100000000000000010000000000010000111111111111001111111111111101111111111111111000111111111111111011111111111011001111111111111001111111111111110000000000000010100000000000000001000000000000011000000000000000011111111111111010111111111111101000000000000001110000000000001110111111111111100100000000000011111111111111111010000000000000000011111111111000000000000000000101111111111111010000000000000000101111111111110010111111111111101100000000000001000000000000000000000000000010100011111111111111000000000000010100111111111111110100000000001001000000000000010100111111111110100011111111110111111111111111111010111111111111110111111111111110100000000000000010111111111111100111111111111110111111111111101011111111111111001111111111111011001111111111111110111111111111100000000000001000100000000000001110111111111111010111111111111110011111111111110110111111111111011111111111111011000000000000010000111111111111101100000000000010110000000000001001111111111111111011111111111111101111111111111100000000000000010011111111111110010000000000000011000000000000111000000000000101010000000000000000111111111110110111111111111101110000000000001001111111111111010111111111111111101111111111110101000000000000100111111111111111111111111111110011000000000000011011111111111110110000000000001011111111111111110111111111111111000000000000000001111111111111010000000000000010000000000000011000111111111111010100000000000001101111111111110100000000000000110000000000000000110000000000001011000000000000010111111111111111110000000000000110000000000000000100000000000000001111111111110011111111111111011111111111111101001111111111101111000000000000110111111111110111110000000000000010000000000000101111111111111111001111111111110010111111111110010000000000000011001111111111110111000000000000000000000000000000011111111111111101000000000000111111111111111101110000000000000001000000000001100111111111111001010000000000000100111111111110011100000000000001011111111111110101111111111111111011111111111111111111111111111101111111111110111000000000000001000000000000100110000000000001101100000000000110011111111111111010111111111110101011111111111111101111111111111101000000000000011100000000000001110000000000000100000000000000101100000000000100110000000000010110000000000001111111111111111110010000000000000000111111111101010111111111111011101111111111100111000000000001001000000000000010010000000000100111111111111111001100000000000100001111111111110000000000000001111011111111111010010000000000000010111111111111010000000000000010011111111111011101111111111110100111111111111111101111111111110101111111111110110000000000000011100000000000010111000000000000111000000000000000011111111111001111000000000000000111111111111111110000000000000000111111111110111100000000000001100000000000001100111111111111110111111111111010011111111111111001000000000000011000000000000011101111111111011011111111111101011111111111111010001111111111110111111111111111101011111111111111111111111111000010111111111111001111111111111010100000000000011100111111111110111011111111111110000000000000101110000000000000000000000000000001010000000000001101000000000001110111111111111111100000000000001110111111111110010111111111111111010000000000010100111111111100011000000000000001101111111111101111111111111111010111111111111101110000000000101010111111111011001111111111110101100000000000001000000000000000100111111111111111110000000000011000000000000001001000000000000001010000000000010100000000000000011100000000000010001111111111011100000000000001001011111111111101011111111111110101000000000000101011111111111111000000000000000000111111111111000011111111111011011111111111110011000000000000001100000000000110010000000000000001111111111111101000000000000100010000000000010010111111111111110111111111111110111111111111110011111111111111011011111111111110000000000000000111111111111110011100000000000011010000000000001001000000000010000000000000000001111111111111110010000000000000010100000000001010000000000000110011000000000001001000000000000000111111111111110111111111111111100000000000000000101111111111101110111111111110001000000000000101111111111111110001111111111111111000000000000001110000000000010111111111111110100011111111111001011111111111101010111111111110110000000000000100111111111111111000000000000000011111111111111111111111111111111011000000000000101011111111110011111111111111010011111111111111110011111111111101001111111111010101000000000000000000000000000010000000000000001101111111111111100100000000000001110000000000000111000000000010010111111111111110001111111111111000000000000001100000000000000101100000000000010000000000000000000000000000000010001111111111101111111111111111010111111111111011110000000000001100000000000001100111111111111111111111111111011110000000000001110100000000000010011111111111111101000000000010000000000000000001111111111111110110000000000000000000000000000111010000000000001000111111111110100011111111111101110000000000011100000000000010011000000000000011001111111111011000111111111111010000000000000000101111111111111110000000000001010111111111110110110000000000000010000000000000110011111111111111110000000000001111111111111111111011111111111111100000000000000100000000000000010000000000000011001111111111111000111111111111010111111111111011001111111111101110000000000000011100000000000001011111111111111111000000000000101100000000000000110000000000000111111111111101100000000000000001111111111111111011111111111110101011111111111101001111111111111010111111111110100111111111111111100000000000010101000000000000001011111111111001111111111111111000111111111110111011111111111111011111111111110110111111111111011000000000000001100000000000000111000000000001000000000000000011110000000000001100111111111111101000000000000001110000000000000101111111111111011011111111111011111111111111101001111111111111011100000000000011011111111111110100111111111111100111111111111011110000000000010000111111111111011111111111111101100000000000011000000000000000111100000000000000111111111111111101000000000000110111111111111110011111111111111001111111111111101111111111111100101111111111110100000000000000010000000000000010001111111111111101000000000001101000000000000101001111111111111000111111111110101111111111110110101111111111111110111111111101111011111111110100101111111111011111000000000000100100000000000000000000000000000100000000000010011111111111111111001111111111110101111111111111101111111111111101110000000000000110000000000001010000000000000000001111111111111001000000000000111100000000001000000000000000000111111111111110011100000000000100110000000000000000111111111111000011111111111001101111111111111100111111111111110111111111111110111111111111110111000000000000010011111111111101111111111111110000000000000010011000000000000011011111111111100101111111111111101100000000000010110000000000001001000000000000000000000000000000001111111111111000111111111111101011111111111110110000000000010001111111111111010111111111111100000000000000001001111111111101111111111111111001001111111111110101111111111110100000000000000000001111111111100110000000000001000011111111111010101111111111110101000000000001000100000000000100000000000000001000000000000000011111111111111110101111111111101010111111111111011111111111111110001111111111011000111111111111111011111111111110011111111111110110000000000001001111111111111011001111111111110010000000000000100100000000000100010000000000010111000000000001001011111111111011011111111111001111111111111111000111111111111111110000000000001111111111111111010000000000001011110000000000000000000000000000100111111111111111110000000000011100000000000001100011111111111111010000000000011101111111111111111111111111111010000000000000000101111111111110111011111111111010101111111111101101111111111111101011111111111111110000000000001010111111111111010000000000000000000000000000100000111111111111010011111111111111010000000000011000000000000000000111111111111101100000000000001010000000000000000100000000000011000000000000000110000000000000100111111111111001000000000000000101000000000000011011111111111110101111111111110110000000000000100000000000000110101111111111101011000000000010001000000000000001011111111111111111111111111111011111111111111101010000000000010001111111111111000011111111111110011111111111110010000000000000101000000000000000000000000000000000111111111111001011111111111010101111111111100111111111111111011111111111111000001111111111100111111111111111001100000000000001000000000000001110111111111110100111111111111110011111111111101001000000000000111111111111111110100000000000001001000000000000010000000000000000100000000000001011000000000000011111111111111010111111111111101011000000000000100100000000000001001111111111111011000000000000010011111111111000011111111111111000000000000001001011111111110110110000000000001000000000000000000000000000000010100000000000011011000000000000001111111111111111100000000000000000000000000000011111111111111110000000000000011101000000000000100111111111111011110000000000011001000000000000010000000000000100011111111111111011111111111111111011111111111111011111111111100011000000000000011111111111111111000000000000000110111111111111011011111111110110111111111111110111000000000001001000000000000110000000000000000000111111111111111011111111111110101111111111100110111111111111011011111111111111010000000000010110111111111111100111111111111110110000000000010101000000000001011100000000000100111111111111110110111111111101100111111111101111100000000000000000111111111111100000000000000010110000000000000010000000000000111100000000000000100000000000001011000000000100001011111111111100101111111111110110000000000011010111111111111100011111111111110101111111111111100011111111111011110000000000000000000000000001000100000000000010111111111111100011000000000000110100000000000001101111111111111100111111111110001111111111110110111111111111101000111111111110001100000000000100010000000000001001111111111111100111111111111111010000000000011010111111111111011000000000000111111111111111110010111111111111000000000000000011010000000000001111000000000001100011111111111111111111111111111010111111111110101011111111111010100000000000011011000000000000001000000000000000110000000000010001111111111111101111111111111110110000000000000010111111111110100111111111110001011111111111001011111111111110100000000000000011100000000000100000000000000000101011111111111111001111111111111110000000000000001100000000000000100000000000010100111111111101000111111111110111001111111111101001111111111111011100000000000001010000000000001111111111111111110111111111111001010000000000001101111111111110110011111111111100110000000000001010111111111110111100000000000101010000000000111110111111111111001011111111110111100000000000000000111111111111010100000000000100010000000001000110111111111110110100000000000011101111111111110100111111111111010011111111110110000000000000000000000000000000010000000000000110100000000000100010000000000000011000000000000011001111111111010110000000000000001011111111111100001111111111001010000000000000011011111111111101010000000000001111111111111110110100000000000011001111111111110101111111111111101011111111111011100000000000001110111111111111100100000000000010100000000001011001000000000001100011111111111010011111111110101001111111111111011011111111110110011111111111001001000000000000000011111111111110101111111111110001111111111111111100000000000000101111111111111101111111111110111011111111111110000000000000000000000000000000101000000000000001100000000000001001111111111111100000000000000110010000000000111000111111111111100111111111111011001111111111101010000000000010011000000000001001110000000000000010000000000001011100000000000000011111111111101100000000000000110000000000000001011111111111111101111111111111011000000000001001110000000000000111000000000000100100000000001011111111111111111110111111111111101000000000000000010000000000010111000000000000010011111111111110100000000000001011000000000000000000000000000110000000000000110000000000000000011111111111110110100000000000000000000000000000011100000000000101000000000000010000111111111111000000000000001101000000000000001100000000000000011011111111111011100000000000000111000000000000100000000000000000100000000000010001000000000001010000000000000001101111111111100000111111111110001100000000000001000000000000000010111111111101001000000000000110001111111111111110111111111111111100000000000001001111111111110011111111111111011100000000000001101111111111101110000000000000111000000000000000001111111111101111111111111111001000000000000101001111111111110001111111111111001011111111111011010000000000000110111111111111111100000000000000000000000001010010111111111101110100000000000100001111111111110100000000000001010100000000000000011111111111011011000000000010000000000000000101111111111111011000000000000000100000000000000000101111111111110101000000000001001111111111111111101111111111110111111111111111001111111111110110000000000000010000111111111101000000000000000010000000000000001100111111111111001000000000000111010000000000011010111111111011100111111111111010000000000000011000111111111111110100000000000001100000000000000000111111111111001011111111111101110000000000001010000000000000010011111111111101011111111111100111111111111111011100000000000011000000000000000110000000000010000000000000000100011111111111110111000000000001110011111111111011111111111111011010111111111111000000000000000000110000000000010011111111111101110111111111110100110000000000000111000000000010011000000000000000001111111111100100000000000000100011111111111111100000000000010100111111111111111011111111111110000000000000000111000000000000000000000000000010001111111111010011111111111110010011111111111100101111111111111100111111111101111011111111111011000000000000010110111111111101111111111111111101110000000000111101111111111110001011111111111000010000000000000111000000000001001011111111111101111111111111001110000000000101101000000000000001110000000000000111000000000000110100000000000000000000000000000001111111111111001000000000000000011111111111111011111111111111010011111111111110101111111111111010000000000000010000000000000110010000000000010110000000000000001100000000000101100000000000010101000000000011111000000000000001110000000001001000111111111111101100000000000011111111111111011101111111111111010100000000000000000000000000011010111111111111101011111111111010100000000000101010111111111101101011111111111101110000000000000000111111111101100111111111111011111111111111111001111111111111110111111111111001101111111111100011000000000001001000000000000010000000000000010110000000000001110011111111111001001111111111111001000000000010100100000000000111100000000000000001000000000000100000000000001000011111111111010001111111111111101100000000000001111111111111111010111111111111111011111111111011101111111111101000111111111110111000000000000000011111111111101110000000000000000111111111111111010000000000001111000000000010101000000000000010110000000000000110111111111110010011111111111110111111111111110000111111111111001000000000001010000000000000001010111111111110011100000000000000110000000000110000000000000000001111111111111101101111111111101101000000000000010011111111111010111111111111110000111111111110100111111111111101000000000000100000111111111110100000000000000000000000000000010111111111111111100000000000000100011111111111110111111111111111111100000000000111001111111111110011111111111110110100000000000000001111111111111110000000000000111011111111111011010000000000011000111111111111100011111111110111010000000000010100000000000000001000000000000011100000000000010000111111111111110100000000000100011111111111111100000000000010100011111111111111011111111110111001000000000000011000000000000011110000000000001010000000000001011100000000000110111111111111110100000000000001011011111111111110101111111111100001111111111111011000000000000000001111111111101001111111111110100100000000000000000000000000001001111111111111101111111111111110001111111111110111000000000001000000000000000000101111111111101111000000000001000100000000000000011111111111110100111111111110010111111111111111000000000000000000111111111110100011111111111011011111111111101110111111111111111111111111111111011111111111110110000000000000001011111111111110111111111111100001000000000000010011111111111111010000000000010100000000000001011000000000000100000000000000101010000000000001011000000000000001111111111111111010111111111111101011111111111001001111111111101111000000000000101100000000000000000000000000100101111111111110111111111111110110000000000000001111111111111101111111111111111101010000000000000111000000000000101100000000000001100000000000101101111111111111100100000000000010111111111111101101000000000001010000000000000001000000000000100010111111111111100000000000001001000000000000101100111111111111101011111111111011101111111111100100000000000010100011111111111110111111111111110011000000000001001011111111111110000000000000000000000000000000001000000000000000001111111111110110000000000001000011111111111111001111111111110101111111111111011000000000000011110000000000000000000000000000000000000000000010010000000000100110111111111101101011111111111101100000000000101010111111111110010000000000000000100000000000011111000000000000000011111111111111011111111111101100000000000000001011111111111100111111111110110110000000000001100000000000000001011111111111010100000000000001000000000000000000001111111111100111111111111111110111111111111010101111111111101000000000000000100000000000000000000000000000000000111111111110011011111111110101110000000000010011111111111110101011111111111111111111111111111101000000000010011100000000000001010000000000010110111111111110110111111111111011010000000000001111000000000001100000000000000110101111111111111010000000000000010100000000000111000000000000001000111111111110001111111111111110001111111111101110111111111111110011111111111011010000000000011101000000000001011011111111111100100000000000010110000000000000001100000000000100111111111111111101000000000000110111111111111010001111111111100000000000000000110011111111111101001111111111110111000000000000100111111111111001111111111111101011000000000000111100000000000001100000000000001011111111111110010100000000000000100000000000101011000000000000000000000000000001110000000000100000111111111111111100000000000001000000000000000111111111111111000000000000000010111111111111111001000000000000000000000000000000111111111111111010000000000000110111111111111110101111111111110111111111111111100000000000000111000000000000001011000000000000101100000000000100000000000000001111111111111111100111111111111001110000000000000111111111111110111111111111111110000000000000000000111111111101001111111111110111011111111111110001111111111101101011111111111010011111111111101000000000000000111000000000000011101111111111101000111111111111000111111111111011110000000000001010000000000001100111111111111110001111111111110011111111111111101100000000001001110000000000011110111111111110101011111111111111011111111111101100111111111111000011111111111111111111111111110110000000000001000111111111111101000000000000000111111111111111011111111111111011110000000000001100000000000010010100000000000001111111111111110100000000000000011000000000000101100000000000001100000000000000111000000000001001000000000000001010000000000000101011111111111011111111111111111110111111111111001011111111111011101111111111110111111111111111100000000000000001000000000000101000000000000000001000000000000100010000000000001110000000000000111111111111111111000000000000000111000000000000010100000000000100111111111111111011111111111111010000000000000011110000000000000011111111111111001100000000000000010000000000100111111111111111011000000000000000111111111111111100000000000000000000000000000011011111111111101001000000000000011111111111111111001111111111111110111111111111100111111111111101111111111111101101111111111111010000000000000011010000000000000000000000000010100100000000000000000000000000000000111111111101100011111111111001111111111111101000111111111110011100000000000010001111111111111101111111111111101100000000010000010000000000011011111111111111100000000000000110110000000000001111111111111110101111111111111000010000000000010110111111111110010011111111111011110000000000101100111111111110100100000000000000111111111111100000111111111111010111111111111101111111111111110111111111111111010100000000000101111111111111010010000000000001100000000000000000001111111111111001000000000000001111111111111110001111111111110010111111111111000100000000000001000000000000000101111111111110000011111111111010110000000000010101111111111111010111111111111111101111111111111010000000000001111000000000000111100000000000000000000000000010111000000000000100101111111111110111000000000000010100000000000110101111111111100100111111111110101100000000000000100000000000010010000000000010011100000000000111010000000000001011111111111111111100000000000000011111111111111010000000000001100011111111111111001111111111100111111111111110011100000000000001011111111111100111000000000000111100000000000101100000000000001111000000000010111000000000001000100000000000011111111111111111000011111111111001111111111111110101111111111111000100000000000010001111111111101010111111111110000111111111111101001111111111110000111111111111101000000000000010011111111111111101000000000000000100000000000100101111111111111101111111111110100111111111111111100000000000000110000000000001001011111111111011001111111111110011111111111110100011111111111100111111111111011101111111111110100100000000000101010000000000110100111111111111110011111111111010011111111111111000111111111110101111111111111000110000000000000101111111111111101100000000000000000000000000100111111111111111100011111111111111000000000000000101000000000000010011111111111111010000000000010001111111111111110000000000000000010000000000000001000000000000011100000000000110100000000000010110000000000000000000000000000100001111111111110100000000000001010100000000000010111111111111110011000000000000010111111111111111101111111111111000000000000000011000000000000011000000000000010000111111111111010011111111111111010000000000000000000000000000100100000000000110000000000000100101000000000000110100000000000110000000000000010001000000000011001100000000000011111111111111101001000000000001010011111111111101110000000000000110000000000000001100000000000000011111111111101011111111111111110011111111111101111111111111100100000000000000010000000000000100011111111111101011000000000000000111111111111111101111111111111100111111111111011111111111111100010000000000000101111111111111100111111111111010111111111111110110111111111101101111111111111100000000000000000011111111111100011111111111111000110000000000010011111111111110100011111111111101111111111111111010111111111111010011111111111110010000000000001100111111111111111100000000000011110000000000110001000000000001011011111111111101101111111111100100111111111101111111111111111111001111111111101111111111111111110011111111111110100000000000000000000000000001011111111111111011001111111111010010000000000001110011111111111100011111111111101101000000000001010100000000000010010000000000001000111111111110000011111111111111001111111111111001000000000010001000000000000101011111111111110111000000000000001111111111111101010000000000010011111111111111110100000000000110110000000000100000000000000001000000000000000000100000000000000000000000000000011111111111111101111111111111110101000000000001001100000000000000001111111111111011111111111111011100000000000000100000000000011011111111111111000011111111111100001111111111111010111111111110010100000000000000011111111111110010000000000000111111111111111010011111111111111101111111111110000000000000000101000000000000000011111111111111010100000000000010100000000000000100000000000000101011111111111110011111111111111001000000000001011000000000000000110000000000000100000000000001000100000000000101010000000000000110111111111111111111111111111100111111111111111111111111111110101111111111111111111111111111111101111111111110010111111111111101110000000000101010000000000000000111111111111011100000000000011101111111111110110111111111111101001111111111101110000000000000100000000000000100001111111111001101000000000000000100000000000111101111111111111100000000000000100100000000000000000000000000001111000000000010000011111111111100111111111111111100000000000001001111111111111110110000000000010000000000000000101111111111110111101111111111101110111111111111101011111111111110000000000000000101000000000000110000000000000000010000000000000111111111111111111011111111111100101111111111101010111111111111000011111111111110000000000000001110111111111111101011111111111110110000000000001000000000000000101100000000000001111111111111110111111111111110111011111111111011111111111111101101111111111111100000000000000100001111111111100010111111111111110000000000000011100000000000000011111111111111100111111111111101110000000000000000000000000000000011111111111101110000000000011000111111111111100011111111111000110000000000000010111111111111111011111111111101000000000000001011111111111111100011111111111101000000000000011100000000000000110111111111111001100000000000010100111111111111101011111111111101110000000000000000000000000000101111111111111101110000000000000000111111111111100100000000000011101111111111111100000000000001100111111111111011010000000000000001111111111111010000000000000010110000000000000111000000000010001100000000000001101111111111111100000000000001010100000000000100000000000000000011000000000000010100000000000010000000000000001010111111111111000111111111111101111111111111101101111111111111100011111111111101101111111111100110111111111111000111111111111011111111111111110001111111111111011000000000000001000000000000001001111111111111111000000000000100100000000000101000111111111111001100000000000000011111111111111000000000000000101011111111111010101111111111111100111111111101110000000000000000001111111111101110000000000000001011111111111110100000000000000110000000000001010111111111111011010000000000000100000000000000111000000000000001001111111111111011111111111111011011111111111101101111111111111000000000000000011100000000000010000000000000010110111111111110101000000000000111000000000000111010111111111111111111111111111000110000000000010000111111111100111000000000000000001111111111110011000000000000101000000000000101001111111111111101111111111111100000000000000001001111111111101011111111111111001000000000000010101111111111110001000000000000110000000000001000101111111111100101111111111111001000000000000001011111111111111101111111111110100011111111111001111111111111110010111111111111000011111111111011110000000000011010111111111101110011111111111110101111111111110010000000000001000000000000000010010000000000000101000000000001001011111111111101001111111111011100111111111110011000000000001011000000000000010010111111111110100000000000000101010000000000011010111111111101000111111111111111111111111111110110000000000000100111111111111100111111111111110100000000000000100100000000001000110000000000100101000000000010000111111111111101011111111111101111111111111111011100000000001100011111111111101110000000000010001011111111110110011111111111101111000000000000011111111111111111100000000000010101111111111110001011111111111100010000000000000111111111111110100011111111111110001111111110110100111111111100110111111111111011000000000000001111000000000000010111111111111101001111111111110011111111111111000000000000000000001111111111110100000000000000011000000000001000011111111111100101111111111111000100000000000011101111111111101001111111111110001011111111110101000000000000101011111111111111010011111111111101110000000000011100000000000001110100000000000001111111111111111000000000000001011111111111111100101111111111111001000000000001001011111111111111101111111111111001111111111111000000000000000100101111111111101110111111111101110111111111111010010000000000000110111111111111001000000000001000111111111111110010111111111101111000000000000111010000000000100010111111111110011000000000000011110000000000100000111111111110000111111111111110000000000000100001000000000000100011111111111111001111111111100101000000000001001011111111111111001111111111111111000000000001011000000000000001111111111111111010111111111111101011111111111101010000000000001111111111111110010100000000001000110000000000011111111111111110010011111111111000100000000000100111000000000001000011111111111100111111111111110000111111111111001011111111111111010000000000100011111111111100100000000000000000110000000000010101000000000011001011111111111111011111111111001100000000000000101111111111111100001111111111111110111111111111010100000000000001101111111111110011111111111110100111111111111101010000000000000010111111111111101100000000000000000000000000010010111111111111101000000000000010100000000000001101000000000000110111111111111111100000000000000101000000000000001111111111111111101111111111101011000000000000011000000000000011101111111111101011000000000000000000000000000000001111111111110101111111111110011100000000000101000000000000000010000000000000111000000000000101111111111111111100000000000000111011111111111110000000000000001010111111111111111011111111111111111111111111110101111111111110111111111111111100111111111111110101111111111111010100000000000100110000000000001111000000000000000000000000000001101111111111101011111111111111110000000000000011010000000000010010000000000000011000000000000100011111111111110000111111111110001000000000000111001111111111111010111111111110100111111111111101110000000000011100000000000000111011111111111111111111111111100010000000000000110011111111111110010000000000001010111111111110111111111111110010101111111111011001111111111111110000000000000001110000000000001100111111111111010100000000001010010000000001001100000000000001001100000000000001011111111111111100000000000000000111111111111101111111111111101111111111111111000011111111111111010000000000001000111111111111011111111111111100111111111111101010000000000001101111111111111101100000000000101111000000000010011000000000000011100000000000101111111111111111110100000000000000001111111111110000000000000001011011111111111100011111111111111001000000000001011100000000000100010000000001000110000000000001100000000000000010001111111111101111000000000000000111111111111111110000000000010011111111111101000000000000000101010000000000011000111111111101111011111111110111001111111111010110000000000000010100000000000000001111111111100111000000000000100100000000000010100000000000000101111111111100110111111111111010111111111111100011000000000000010100000000000010001111111111010110000000000001001011111111111111100000000000000101000000000000101100000000000100110000000000101100111111111111111111111111110101101111111111111101111111111111011011111111100110111111111111000111000000000000001000000000000001110000000000100000000000000001001000000000000011000000000000010010111111111111010111111111111001110000000000000011111111111110011111111111110101001111111111010101000000000000000111111111111011101111111111111001000000000010111100000000001100000000000000111011000000000000001000000000000000000000000000011111000000000000111011111111111101110000000000000001000000000000000011111111110111110000000000000000000000000000011011111111111111101111111111110100000000000000000100000000000000000000000000100000111111111100101100000000000000010000000000100111000000000000111011111111111101100000000000001010111111111111111111111111111100111111111111101111111111111111101011111111111100000000000000001111111111111101101111111111111010011111111111101001111111111111001100000000000010000000000000000011111111111110101100000000000000101111111111111111111111111100010011111111110110101111111111000110111111111110010100000000000010100000000000010111000000000001111100000000001001100000000001001000111111111101011100000000000010010000000000000100000000000001101111111111111110110000000000010101000000000001110100000000000011010000000000001010111111111101000011111111111001001111111111001100000000000000011000000000000010000000000000001001000000000001010000000000000010000000000000000100000000000001001111111111111110000000000000000111000000000001010111111111111101111111111111111111000000000001001111111111111110100000000000100100000000000001110100000000000011100000000000010011000000000001101111111111111110001111111111110110000000000000111111111111110101111111111111101100111111111100100011111111111011111111111111100011000000000000000111111111111010101111111111111010111111111111110100000000000000010000000001001100000000000000000111111111110000001111111111011000111111111110001011111111110111010000000000000011111111111101100100000000000101010000000000110000111111111111010100000000000110101111111111011111000000000000110111111111111011111111111111111110111111111110100000000000000001101111111111100101111111111100111111111111111011111111111111100101111111111110110111111111111010101111111111111001111111111111011100000000000011010000000000001001111111111111100111111111111001101111111111110101000000000000110100000000001001001111111111110010000000000001111000000000000001010000000000100101000000000010110000000000000111110000000000010101000000000001101000000000000111100000000000010100000000000000010100000000000011110000000000011010111111111110111100000000000000001111111111101111000000000000000000000000000100011111111111101110111111111111001111111111111010101111111111111100111111111110000011111111111100000000000000000110111111111110001000000000000001010000000000011100000000000011000000000000000010100000000000000111111111111101100111111111111111001111111111100011000000000000010111111111111011110000000000010100111111111111100000000000000000110000000000101011000000000000001000000000000010100000000000011010000000000000110111111111111101010000000000010101111111111111110000000000001010100000000000001000111111111110111011111111111110001111111111010110000000000001100100000000000011110000000000011010111111111111001111111111111000000000000000010011111111111110101111111111111001101111111111001010111111111111001111111111111110010000000000100111000000000001010100000000000011000000000000011110000000000001101000000000000010101111111111110111000000000000100111111111111111101111111111101011111111111110110111111111111111111111111111110100000000000000010100000000000011100000000000000011111111111111001100000000000010011111111111111000111111111110111000000000000000111111111111110111000000000000100100000000000100101111111111101110000000000001000100000000000011111111111111111111000000000001001000000000000001101111111111111101000000000000011111111111111010101111111111110010111111111110011011111111111011111111111111111100000000000001010011111111111010110000000000000000000000000001000100000000000010110000000000010001000000000000111111111111111111110000000000001101111111111111100000000000000001010000000000010110000000000010110100000000000001110000000000010110000000000001010111111111111111011111111111101111111111111111111011111111110110111111111111101110000000000000010011111111111101001111111111111000111111111111111011111111111101111111111111110011000000000000001100000000000010000000000000001111111111111101010011111111101110001111111111000100111111111101100100000000000010101111111111111101111111111111100011111111111111000000000000111011111111111111010100000000000000000000000000011111000000000000100100000000000100001111111111101110000000000001100011111111111110011111111111010011111111111101001111111111111101101111111111110111000000000000100000000000000000010000000000110010000000000000100011111111111100011111111111110000000000000000000011111111111101011111111111111110000000000001010100000000000010000000000000000010000000000000011011111111111011010000000000000100000000000000110100000000000100000000000000000000111111111111101111111111111111101111111111111110000000000000001011111111111100011111111111101101111111111111111100000000001000001111111111111111111111111110011100000000000001001111111111111010000000000001101111111111111000111111111111111111000000000000110011111111111111000000000000001010111111111111000011111111111001111111111111100001111111111111000100000000000000010000000000000100111111111111001011111111111110001111111111101010111111111111110111111111111111011111111111100001000000000001111000000000000001010000000000010100000000000001000011111111111011001111111111110001000000000000001011111111111111011111111111101111111111111111000111111111111101001111111111110100111111111111010011111111111111011111111111111110000000000000100000000000000000010000000000000110000000000001101000000000000010100000000000110000000000000010110100000000000111010000000000001001000000000001100111111111111011000000000000001001111111111111101111111111111101100000000000001100111111111111001000000000000000010000000000001000111111111111011011111111111101100000000000000111000000000000010100000000000000011111111111111101111111111110110111111111111110101111111111010011111111111111111011111111111101101111111111111001111111111111010100000000000001110000000000001000111111111111110100000000000000010000000000000000000000000000100011111111111101100000000000000000111111111111011011111111111111101111111111110101000000000000010100000000000100010000000000000001111111111111000111111111111100111111111111111100111111111111110100000000000000100000000000010011000000000001111111111111111011100000000000001110111111111111011011111111111100100000000000000010000000000000000000000000000100010000000000001001000000000000100000000000000011011111111111111010111111111111101100000000000000100000000000000001111111111111000011111111111111100000000000001100111111111110111100000000000000000000000000000100111111111111101100000000000001100000000000000000000000000000010111111111111110111111111111110100000000000000110011111111111111110000000000000000000000000001000111111111111110100000000000000010111111111111001000000000000001011111111111110100000000000000010100000000000001000000000000100010111111111111110000000000000000100000000000000111000000000000011111111111111101111111111111100100111111111110111111111111111110011111111111011010111111111111001011111111111101001111111111111011111111111111011111111111111110101111111111110100000000000000011111111111111111000000000000001111000000000000000111111111111010101111111111111110111111111111001111111111111110100000000000010011111111111110111111111111111100111111111111011110111111111111100000000000000011000000000000000000000000000000000000000000000000011111111111101101111111111111001011111111111100110000000000001110000000000000010011111111111110010000000000000000000000000000000000000000000001010000000000010011000000000000110000000000001101001111111111111001000000000000000100000000000001111111111111110100000000000000011011111111111101001111111111111010111111111110111100000000000001110000000000001100000000000000001011111111111001001111111111110101111111111111110111111111111100101111111111110010000000000000001000000000000010100000000000000100111111111111100000000000000011010000000000001111000000000000000100000000000011100000000000100100000000000000010000000000000000010000000000001101111111111111101000000000000001011111111111111001000000000000100100000000000000011111111111111010111111111111111111111111111100110000000000000001000000000000001011111111111010111111111111101110111111111110101111111111111101011111111111111000000000000000100100000000000001001111111111110010111111111110101111111111111111001111111111111011000000000000011111111111111110100000000000001011111111111111111100000000000010011111111111110011111111111111111011111111111111010000000000001110111111111110111011111111111111110000000000000000000000000000000100000000000001110000000000001111111111111111111011111111111100011111111111101110111111111111101000000000000011110000000000000001111111111110101111111111111111001111111111111001000000000000011000000000000010001111111111111100000000000000010111111111111110110000000000010010000000000000100011111111111101000000000000011001000000000000000011111111111110100000000000010100111111111111001111111111111101110000000000001010111111111111000111111111111101000000000000001001111111111111001011111111111011110000000000000001111111111110111111111111111111101111111111111101111111111111001100000000000010010000000000010101000000000000100011111111111111001111111111110100000000000000110100000000000001011111111111111110000000000000001000000000000110100000000000011011111111111111011100000000000011100000000000011001000000000000110000000000000001110000000000000000000000000000011011111111111010111111111111111010000000000000001111111111111111001111111111111111000000000000100011111111111011101111111111111110000000000000111100000000000100011111111111111001111111111111101111111111111110110000000000011000111111111110111000000000000000111111111111111010111111111111100011111111111010111111111111100101111111111111100011111111111110001111111111110101111111111111111011111111111111110000000000000010000000000001000011111111111100101111111111101100000000000001000111111111111111001111111111100001111111111110100100000000000001010000000000010100000000000001011011111111111101000000000000000101000000000001010111111111111111100000000000001001000000000000000111111111111110011111111111100111111111111111101100000000000001100000000000000011111111111111111111111111111101101111111111101111111111111111101100000000000000000000000000000001000000000000001011111111111100101111111111011100000000000000011100000000000011110000000000000000000000000001000000000000000000010000000000000111111111111111010100000000000001010000000000000011111111111111001011111111111111100000000000001101000000000000110000000000000001001111111111111111000000000001100100000000001011000000000000100110000000000000110100000000000011101111111111111111000000000001001100000000000000100000000000000010000000000000000011111111111011001111111111111100000000000001001000000000000000100000000000000101111111111111101111111111111101011111111111111110111111111111011100000000000001101111111111111101000000000000011000000000000001010000000000001110000000000000011000000000000011000000000000001010000000000000000011111111111110111111111111101010111111111111010011111111111100100000000000001011111111111110000011111111111001101111111111111110000000000000010100000000000010110000000000001011000000000000100011111111111001100000000000000000000000000001001011111111111111010000000000001001000000000000100111111111111110111111111111111110000000000000001111111111111111100000000000001110000000000000011100000000000110111111111111100000111111111111110000000000000001101111111111111111000000000000001000000000000000100000000000000000000000000000000000000000000000000000000000000111111111111111011100000000000110010000000000011101111111111111110100000000000000001111111111111101111111111101101011111111111101000000000000000100000000000000001000000000000110110000000000000101111111111110110100000000000000000000000000001100000000000000001011111111111101101111111111111100111111111111110100000000000001010000000000000101111111111111111000000000000001110000000000010011000000000000000011111111111111000000000000000110111111111111101011111111111100111111111111011110111111111111101100000000000000001111111111101111000000000000011011111111111101010000000000010000111111111111010011111111111111001111111111111000111111111111101011111111111100011111111111111100000000000000010111111111111111110000000000000110000000000000111011111111111101001111111111111100000000000000100111111111111110001111111111111110000000000000010000000000000011111111111111101111000000000000010100000000000000000000000000001010111111111111101000000000000000011111111111110101000000000000010011111111111100111111111111100001000000000001000100000000000110010000000000010010000000000001001011111111111111101111111111111111000000000000111000000000000001110000000000000000111111111111011100000000000011100000000000010101000000000001001000000000000011010000000000000010111111111101110011111111111101011111111111111110111111111111111111111111111100111111111111100101000000000000000000000000000000001111111111101001000000000000011000000000000010101111111111100111000000000001010100000000000011000000000000001000000000000000011100000000000000101111111111111000111111111111100111111111111110000000000000000111111111111110101111111111110001111111111111010001000000000001111111111111111100001111111111110111111111111111011000000000000011110000000000010000111111111111001011111111110100111111111111111011111111111111000100000000000010011111111111101010000000000010111100000000001011100000000000000011111111111110100011111111111001001111111111011100111111111111010011111111111101100000000000000010000000000000000000000000000000110000000000100110000000000000000000000000000011110000000000000010000000000000010100000000000000001111111111110010111111111110001111111111111111001111111111110111111111111111100111111111111100011111111111101010111111111111001000000000000111101111111111110011111111111011011000000000000111110000000000101011000000000001100111111111111001101111111111111101111111111111001100000000000010101111111111100000000000000001010011111111111111111111111111101100000000000000100000000000001001100000000000001111111111111101111000000000000001101111111111100000111111111111000111111111111100001111111111101110111111111111111111111111111100011111111111101110000000000000001111111111111100010000000000101011000000000010000100000000000001111111111111110111111111111110111100000000000010101111111111100101111111111110011000000000000010001111111111111101000000000010011000000000000010001111111111100100111111111110000011111111110101101111111111110000111111111111001011111111111111110000000000000000000000000001101000000000000110111111111111111110111111111111010000000000000000101111111111111011000000000000010011111111111101110000000000000001111111111101110111111111110001110000000000001010111111111101101011111111111011111111111111010110111111111111001100000000000001111111111111100111000000000001100100000000000110010000000000100001000000000000001011111111111101011111111111101111111111111111111100000000000000011111111111111000111111111111110011111111111100000000000000001101000000000000110100000000000111110000000000000001000000000000011011111111111010111111111111111100000000000011100000000000000001111111111111111001111111111111011100000000000010010000000000100011111111111111101000000000000000010000000000000000111111111111101111111111111010101111111111011011111111111111011111111111111010111111111111101101111111111111010011111111111110110000000000011011000000000000100000000000000000101111111111101001111111111110001111111111110101011111111111100100000000000001101111111111111110001111111111110101111111111111000100000000000001000000000000000011111111111111001011111111110110111111111111101110111111111111100011111111111011001111111111011110111111111111101111111111111101111111111111100000111111111111011000000000000010101111111111110001111111111111111111111111111101001111111111110101000000000000100100000000001101100000000000010011000000000000101000000000000100000000000000101010000000000000111011111111111101000000000000010111111111111110011000000000000110000000000000010110111111111101110000000000000001011111111111100000111111111111010100000000000000000000000000000100111111111111000100000000000010101111111111110101000000000000000100000000000111110000000000001101000000000000000100000000000101011111111111110000000000000000011111111111111110111111111111000000000000000000100111111111111010011111111111101101000000000010000011111111111100000000000000010001000000000001000100000000000000101111111111110000111111111111111100000000000110010000000000111001111111111111001100000000000110110000000000000110111111111100110000000000000000001111111111111011111111111111001100000000000110100000000000010011000000000000000000000000000010000000000000000000111111111110000111111111111010011111111111101101111111111110100111111111111101001111111111101010000000000000110011111111111101110000000000010001000000000000011100000000000011011111111111100000000000000010000111111111111111011111111111111010000000000000110011111111111011100000000000001100000000000001001000000000000010001111111111111100000000000000000011111111111101101111111111111101111111111111100011111111111110110000000000000000111111111111100000000000000010010000000000001011000000000010111000000000000100001111111111111000111111111111111111111111111100100000000000100001111111111101011011111111110100100000000000010101000000000001011111111111111111100000000000000110000000000000110100000000000000011111111111101010000000000000111011111111111111111111111111111000111111111111101100000000000001001111111111110001111111111111111011111111111111100000000000000000111111111101110111111111111110101111111111111001000000000000101011111111111100010000000000000101111111111101000100000000000010100000000000001001111111111111111000000000000000101111111111111111000000000001111000000000000100111111111111110011000000000001001000000000000000111111111111100000000000000000011011111111111101100000000000001010000000000000111100000000000010101111111111100100000000000000010000000000000010001111111111011110000000000010110000000000001000000000000000000110000000000001100000000000000010101111111111101000000000000001111100000000000000010000000000001001111111111110000111111111110101001111111111110000000000000001001000000000000100111111111111010001000000000010110011111111111110111111111111100101111111111111010111111111110011011111111111101100111111111111101111111111111111111111111111111010000000000001111100000000000010100000000000000010111111111111111111111111111110000000000000001000000000000000111011111111111110000000000000001010111111111111111011111111111111111111111111101110000000000000000100000000000000001111111111101010111111111111110000000000000011101111111111110000000000000001011000000000000001000000000000000100000000000000000100000000000000100000000000001001111111111101110100000000000100011111111111111011000000000000000011111111111111101111111111100100111111111111000100000000000100100000000000100000000000000000101000000000000100110000000001000011111111111101111000000000000011010000000000001010000000000000000011111111110100011111111111001101111111111111011111111111111100111111111111111011111111111111010111111111111111010000000000001100111111111110101000000000000001100000000000000111000000000010110100000000000011111111111111010101000000000010011100000000000101111111111111111001000000000000100111111111111110110000000000010000000000000001001100000000000100110000000000010111111111111111101100000000000001000000000000000011000000000000000011111111110110110000000000000010111111111111001011111111111110111111111111111001000000000000101100000000000000100000000000010000111111111111111011111111111111010000000000001111000000000001111000000000000000001111111111111100111111111110111100000000000100101111111111111011000000000000010111111111111010111111111111111100111111111110100111111111110111001111111111111011111111111111100100000000000000011111111111111100111111111111101100000000001000100000000000000111111111111111110100000000000000100000000000010010111111111110100100000000000010100000000000011011000000000000001100000000000000101111111111111111000000000000000011111111111111110000000000100011111111111111111000000000000010111111111111111001000000000000100000000000000101011111111111101100111111111111111000000000000100000000000000001101000000000000011011111111111011000000000000100001111111111101100011111111110110101111111111111110111111111111010111111111111110000000000000001001000000000000101011111111111110000000000000000101111111111111101100000000000001011111111111010100111111111111010011111111111110110000000000001101000000000000110011111111111111101111111111111110000000000000000000000000000000100000000000001011000000000000011000000000000001001111111111111111111111111111100111111111111010111111111111110000111111111110111011111111111100111111111111110011000000000000000000000000000010111111111111110000000000000000101100000000000101101111111111110101000000000000010011111111111110010000000000000100111111111110111111111111111011000000000000000100111111111111010100000000000010111111111111111010111111111110100011111111111100000000000000000110000000000000011011111111111001001111111111111101111111111110111011111111111101110000000000000000000000000000110100000000000000101111111111111011000000000001010111111111111101101111111111111000111111111111100011111111111101010000000000001111000000000001100000000000000101110000000000011010000000000000100011111111111011101111111111101111000000000000100111111111111111011111111111111010000000000000010100000000000001101111111111101010000000000010001011111111111100111111111111110101000000000000010111111111111110110000000000000000000000000000101100000000000110100000000000001010000000000000110100000000000011101111111111111011000000000000111100000000000000111111111111101000111111111110000011111111111010101111111111111101111111111111010000000000000000010000000000000010000000000000111011111111111110001111111111110111111111111111110000000000000000001111111111111111000000000000010100000000000001111111111111101100000000000001000011111111111110000000000000000011111111111111011111111111111011000000000000000111000000000000000100000000000000001111111111100101111111111111010100000000000001111111111111111110111111111111011100000000000000110000000000000101111111111100110000000000001000100000000000001111111111111110101111111111111111000000000000001100000000000010001000000000000011100000000000001111111111111111101000000000000010100000000000110000111111111111110000000000000001011111111111111100111111111111011111111111111010011111111111010101111111111111001011111111111001011111111111110001111111111111001111111111111110011111111111111011000000000000001100000000000000110000000000001110000000000001011011111111111101001111111111101100000000000010011000000000000100000000000000000011000000000000001000000000000000110000000000000010000000000000110111111111111110111111111111111010111111111110011011111111111100001111111111111001000000000000000011111111111110110000000000001001000000000001100011111111110011111111111111101101000000000001010100000000000000001111111111100000111111111111000111111111111111011111111111111110111111111111001000000000000000001111111110111111000000000011001111111111110110110000000000000000000000000010110000000000000111010000000000011110000000000000101111111111111101110000000000011100000000000010110000000000000111000000000000010001000000000000011011111111111011010000000000100001000000000001100000000000001000010000000000101010000000000010101111111111111010111111111111101001000000000000010100000000000001000000000000000111000000000010001100000000000001101111111111110101000000000010000011111111111111100000000000010001000000000000011111111111111101111111111111111001000000000000000000000000000111011111111111101100000000000001000111111111111101000000000000000001111111111110101000000000000101100000000000010010111111111101110111111111111011011111111111101001111111111111011111111111111011111111111111011111000000000000100000000000000100010000000000000110111111111110011100000000001010000000000000100101111111111111010100000000000000001111111111111100111111111111001011111111111100110000000000011001111111111101011111111111110111000000000000111100111111111110101100000000000011100000000000000011111111111101111011111111111101011111111111011101111111111110100111111111111011111111111111110100111111111111011000000000000101101111111111110010000000000010000000000000000110001111111111101101000000000000000011111111111111001111111111101000111111111111111111111111111001101111111111111000000000000000000111111111110101101111111111110010000000000011000100000000001010100000000000011011000000000001110100000000000000010000000000001010111111111110110111111111111110011111111111010011111111111110010011111111110001000000000000010110111111111110100000000000000011110000000000100001000000000010010100000000000010001111111111100100000000000001111000000000000011111111111111111011111111111111010000000000000011111111111111101111000000000000001011111111111100011111111111101100111111111110001011111111110100110000000000101010111111111110001011111111111101100000000000011110111111111111001011111111111011011111111111100101111111111101110111111111111100110000000001001000111111111110101011111111111101101111111111110011000000000000000011111111111011100000000000010001000000000000000111111111111110100000000000101010000000000000000111111111111011111111111111111110000000000000010111111111111111110000000000010001111111111111011011111111111000001111111111100111000000000001100100000000000111010000000000001111000000000011101100000000000011101111111111111111000000000001001011111111111101001111111111111001000000000001110100000000000000011111111111111110000000000000111011111111110101101111111111100110111111111111011011111111111010111111111111011010111111111111101111111111111100001111111111100111000000000001100000000000001001000000000000011010111111111111010011111111111110110000000000011000000000000000100011111111111001001111111111111111111111111111100011111111111110111111111111100110000000000001110011111111111100110000000000001111111111111111111111111111111110011111111111101011000000000000111111111111111011000000000000011001000000000001011111111111110111110000000000111111111111111110111000000000000011010000000000000101000000000001101000000000000000011111111111110010111111111110001111111111111111100000000000101111111111111101001100000000000000000000000000011101111111111111101011111111111010111111111111100101111111111110101100000000000000100000000000100110000000000000011011111111111000111111111111111100111111111110111000000000000111000000000000010010111111111110001000000000000010100000000000010110111111111111011000000000000010100000000000000111000000000001001000000000000100000000000000001101111111111111101000000000000111101111111111101111000000000000110011111111111111010000000000001001000000000000110111111111111100100000000000000010000000000011100000000000000101111111111111011101000000000001100011111111111011011111111111111101111111111111011011111111111111101111111111101010000000000000101111111111111011001111111111100011111111111111100011111111111101011111111111100101000000000001011011111111111101111111111111111010111111111110010100000000000001101111111111100010000000000000000000000000000001001111111111110010000000000011011000000000000000101111111111110110000000000001101100000000000101110000000000011010111111111111110100000000000111110000000000000111111111111111100000000000000000111111111111110010111111111111000111111111111111000000000000000001000000000000101111111111111100010000000000010010000000000000110000000000000001000000000000001010000000000001010011111111111101101111111111011100000000000000010111111111111111011111111111100001000000000010111100000000000001001111111111110100000000000000011011111111111111100000000000111000000000000000001111111111111011011111111111101101111111111111111011111111111110100000000000001010000000000000011000000000000011010000000000010100000000000011001011111111111111110000000000001010111111111110111111111111111101010000000000100101000000000010001100000000000000111111111111110010000000000000101111111111111010101111111111001100111111111110001011111111110100101111111111010111000000000000111011111111111110011111111111101000000000000001001011111111111010101111111111101100000000000000101100000000000000100000000000011110111111111110010100000000000001001111111111100101000000000000010011111111111100110000000000011100111111111110111000000000000011100000000000100110000000000000010000000000000101100000000000011010000000000001110011111111111110001111111111011011000000000010011100000000000101011111111111100101000000000000110011111111111110000000000000011011000000000001010100000000000000001111111111111101000000000000000100000000000001101111111111111101000000000001000011111111111110100000000000000001000000000001010011111111111010111111111111111111000000000001100000000000000011111111111111101111111111111110110100000000000001010000000000011110111111111111001011111111111111011111111111111110111111111110101011111111111001110000000000100001111111111100111100000000000000001111111111111111000000000000101000000000000010011111111111111110000000000001011111111111111110100000000000100000111111111111001111111111111101100000000000010011111111111110110111111111111001001111111111111110111111111101111111111111111010110000000000000011111111111111010100000000000110011111111111000100111111111110111011111111111101011111111111111010111111111111011011111111111110001111111111101111111111111111001011111111111110111111111111111110111111111111010011111111111101111111111111111011111111111110111000000000000000000000000000101100000000000000100100000000000010100000000000100110000000000010000100000000000010110000000000000110000000000011010000000000000101001111111111100100000000000000010000000000000001011111111111110001000000000001010100000000000100001111111111010001000000000001010011111111111011001111111111100000000000000001000011111111111110101111111111101011111111111111101011111111111111001111111111110000000000000000101111111111111101000000000000000000000000000001001011111111111100101111111111110101111111111111111111111111111101010000000000010011111111111111011100000000000100111111111111110011111111111110001011111111111000010000000000011011111111111110111100000000000010100000000000010010000000000000001000000000000010000000000000000000000000000001011000000000000100110000000000000010000000000001111100000000000110000000000000001110000000000000011111111111111000000000000000000000000000000011111100000000000010000000000000011101000000000000110100000000000000111111111111111100111111111111111100000000000100000000000000000100111111111110000011111111111101100000000000001110000000000001010111111111111101000000000000001111111111111111101111111111111011010000000000010011111111111111101100000000000000100000000000000100000000000000000111111111111110010000000000000101000000000001101100000000000010001111111111110101111111111110001011111111111000000000000000010011000000000000101011111111111110011111111111110110111111111111011000000000000000000000000000010111111111111111100011111111111011100000000000000011111111111110101100000000000010001111111111111100111111111101111111111111111011010000000000010011111111111111111011111111111110101111111111111011000000000001100111111111111101010000000000011100111111111111100100000000000000101111111111111010111111111010101011111111111000110000000000000000111111111111110011111111111110101111111111110010111111111111111011111111111100011111111111101010000000000000000000000000000110010000000000000011000000000001111000000000000101111111111111111010000000000000000000000000000100100000000000011110111111111110010011111111111100001111111111110001111111111111111011111111111101110000000000010011000000000000101000000000000111000000000000001100000000000010001100000000000111011111111111110100111111111111010000000000000110100000000000011010111111111111010100000000000011111111111111111000111111111110010011111111110110001111111111111111111111111110101011111111111100111111111111101011000000000000000011111111111110100000000000000101111111111100111111111111111001000000000000001111111111111101101000000000000000100000000000001101000000000000100100000000000011001111111111101111000000000001000111111111111010100000000000001011000000000000011011111111111101011111111111110000111111111111001100000000000010010000000000000000111111111111001100000000000010100000000000100010000000000010010000000000000010010000000000001101000000000001011000000000000010001111111111110101000000000001110100000000001101110000000000000000111111111111010000000000000101101111111111110010111111111111111011111111111110101111111111101010000000000001110100000000000010110000000000000000000000000001011000000000000000000000000000001010111111111111011100000000000000000000000000000101111111111101110111111111111000110000000000001011000000000000001000000000000011100000000000000000111111111110011011111111111110000000000000000111000000000000000000000000000101111111111111111111000000000000111100000000000110011111111111111110000000000000010000000000001000001111111111111110111111111101111011111111111111100000000000101010111111111110001111111111111110100000000000000011111111111110101111111111111111000000000000100000111111111101010100000000000000010000000000000111000000000000100000000000000110001111111111111011111111111111000000000000000101100000000000011101111111111111011000000000000010111111111111110111000000000000000011111111111101100000000000001000000000000000010100000000000010110000000000000110111111111110100111111111111011101111111111100111000000000000011000000000000000111111111111111101111111111111110011111111111000011111111111111000000000000000111011111111111010110000000000000101111111111111010111111111111010011111111111110101000000000000111011111111111111101111111111110001000000000000000000000000000001001111111111111111000000000000011000000000000110010000000000000011000000000000110011111111111100001111111111100101000000000000101100000000000000000000000000010100111111111111011111111111111111100000000000000110111111111110101111111111111101011111111111111101000000000000100100000000000110011111111111111111000000000000101000000000000010010000000000001111111111111111100111111111111011111111111111110011111111111111011000000000000001011111111111111010000000000000000011111111111110000000000000011001000000000001011100000000000000100000000000100000000000000001001011111111111111110000000000001010000000000000110000000000000011000000000000001101111111111111111100000000000100011111111111111110111111111111110000000000000100110000000000010010111111111111111000000000000100110000000000010001111111111111011000000000000000001111111111100001000000000000011111111111111111001111111111101100000000000000101111111111111010100000000000000000111111111111101111111111111111000000000000001000111111111111001011111111111011111111111111111011000000000000010100000000000000001111111111111101000000000000110011111111111101101111111111110100111111111110010011111111111110011111111111101001000000000001000011111111111111001111111111101101000000000000001011111111111100001111111111111001111111111111001111111111110111000000000000100010111111111111110111111111111110010000000000000000111111111111110100000000000001010000000000010001000000000000110000000000000001101111111111111010111111111110011111111111111101011111111111111100000000000001000011111111111101001111111111110010000000000001011111111111111100011111111111101100000000000000101111111111111111011111111111111111000000000000000000000000000000000000000000001010111111111110100100000000000011000000000000011111000000000000101111111111111110111111111111111110111111111111011000000000000010001111111111101011000000000001000011111111111110110000000000001100111111111110111000000000000011001111111111101111111111111111100111111111111111010000000000000001111111111110011100000000000010011111111111111110000000000000001000000000000000010000000000000010111111111111000011111111111100001111111111110001000000000001111111111111111111111111111111110110111111111111001011111111111110010000000000001001111111111111101111111111111110011111111111110010111111111101110100000000000011010000000000010011111111111110011000000000000000101111111111111000111111111111110100000000000001000000000000000000111111111110110100000000000100000000000000100010000000000000101000000000000011010000000000001111000000000000011100000000000010000000000000000001000000000000000000000000000011100000000000000111111111111110011011111111111111110000000000010100111111111111101011111111111101110000000000001111000000000000110111111111111101101111111111111000000000000000100111111111111011111111111111111111000000000000100111111111111101101111111111110101000000000000001111111111111010111111111111111010111111111111100100000000000011001111111111110110000000000000100100000000000010001111111111111010111111111111101111111111111010111111111111100100111111111111001100000000000001000000000000000000000000000000101000000000000010101111111111111100111111111111100011111111111100001111111111111110111111111110111100000000000010010000000000000011000000000000000000000000000001010000000000000001111111111111111000000000000010100000000000101010111111111110100100000000000010110000000000000011111111111111101011111111111111010000000000001110111111111110100011111111111011100000000000001001000000000000001000000000000001000000000000000000111111111111100100000000000000010000000000001000111111111110001100000000001010110000000000000110111111111111110100000000000010000000000000001101111111111111001000000000000011111111111111111001000000000000101011111111111101110000000000000100111111111111011000000000000000111111111111111000000000000001100100000000001000010000000000011110000000000000010011111111111111001111111111110011111111111111101000000000000011111111111111111111111111111101011100000000000100001111111111111010000000000001001100000000000010001111111111111110000000000000011111111111111101000000000000000100000000000000101000000000000100011111111111111111111111111110111111111111111100110000000000001011111111111111001011111111111100010000000000000000111111111111101011111111111011101111111111110111111111111110100100000000000010100000000000010111111111111101101000000000000000100000000000000010000000000000001000000000000111001111111111111010000000000011001011111111111001100000000000000100000000000001100000000000000010010000000000000010000000000010100111111111111111010000000000010001111111111110100100000000000101100000000000001010111111111111011011111111111110010000000000011000111111111110100011111111111101001111111111100001111111111110110100000000000011100000000001000000000000000000000011111111111110000000000000010001111111111111011111111111111111000000000000001001111111111101111100000000000011110000000000111000111111111110011000000000000000000000000000001000111111111011110000000000000010010000000000001011000000000000001000000000000100111111111111110110111111111111000011111111111101110000000000001101111111111111110011111111111111011111111111100011000000000000000000000000000111001111111111111101111111111111011011111111111011000000000000000011111111111111110111111111111100111111111111111010000000000000111000000000000010011111111111111111000000000000001011111111111111100000000000000000000000000000001100000000000000001111111111111101000000000001000111111111111011001111111111110001111111111101110100000000000110000000000000000001000000000000111100000000001001010000000000010100000000000000100111111111111000101111111111101100000000000001011011111111111100100000000000001100111111111110101000000000000001010000000000010010111111111111011011111111111100010000000000100001000000000000010100000000000100100000000000001101111111111111011100000000000100001111111111111101000000000001101000000000001001010000000000011100111111111111011011111111111000111111111111110011000000000011000100000000000110110000000000000000000000000000111000000000000000010000000000000111000000000000100011111111111101101111111111110011111111111111100000000000000001110000000000000011111111111110011100000000000100111111111111100001111111111111100000000000000000110000000000000001111111111110011100000000000000001111111111110111000000000000000000000000000010101111111111110001111111111111111011111111111111100000000000010000111111111111110000000000000010111111111111101110111111111110011100000000000001001111111111111100000000000000100011111111111101111111111111100000111111111111010011111111111101011111111111111011111111111111001000000000000010111111111111100110111111111110110100000000000001110000000000000101000000000000011100000000000000011111111111110110111111111101000011111111111011000000000000000011000000000000111100000000000000010000000000101000111111111111110111111111111001101111111111111001000000000001101000000000000010000000000000000000111111111110111011111111111111100000000000000010000000000010101000000000000100000000000000000110000000000010000100000000000100010000000000001000111111111111111011111111111011101111111111100101000000000000111100000000000001010000000000001001000000000000110000000000000011111111111111101011111111111110111011111111110101001111111111101101000000000001111111111111111110100000000000001100111111111111010011111111111110010000000000011111111111111111101011111111111110001111111111000110111111111110101100000000000000010000000000001111111111111111011000000000000001000000000000101011111111111111100100000000000000110000000000000001000000000000010000000000000011010000000000000000000000000000011111111111111001101111111111011010000000000000000011111111111111010000000000010110111111111111001011111111111101100000000000001011111111111111010011111111111101110000000000010110000000000000001011111111111101000000000000000101111111111111000100000000000000111111111111111000111111111100101111111111111100101111111111110101111111111111011011111111111110000000000000001100111111111111010111111111111100101111111111111010000000000001011011111111111101000000000000010111000000000001111100000000000101000000000000100001111111111111001000000000000010100000000000010110111111111110100111111111111100101111111111110101111111111111111000000000000001010000000000101001111111111110000111111111111011101111111111010011000000000000010000000000000000100000000000010000111111111111111000000000000101010000000000010010111111111101101111111111111100101111111111100100000000000000001011111111111011010000000000100110111111111110100011111111111110111111111111111011111111111110011100000000000001100000000000000110111111111101111011111111111110100000000000000000111111111111011000000000000000001111111111111110000000000001010100000000000000001111111111111010000000000000010000000000000001010000000000010100000000000000010111111111111110111111111111101110000000000001000011111111111111101111111111111001111111111110001011111111111101000000000000010000000000000000000111111111111110101111111111111111000000000000111100000000000010011111111111101010111111111111111100000000000110011111111111110011000000000001001111111111111110111111111111110110000000000000000111111111111101110000000000000001000000000010101011111111111101111111111111101011000000000001010100000000000001100000000000001010000000000010000111111111111111100000000000000000111111111101010011111111111100011111111111110000000000000001001111111111111100001111111111111101111111111111110100000000000011000000000000101011000000000001111011111111111011111111111111110101000000000000010000000000000100000000000000001111111111111111011111111111111111000000000000001110111111111110011100000000000001100000000000101101111111111111100000000000000001111111111111110111111111111110101011111111111101011111111111100011111111111111110011111111111101100000000000000001111111111111001100000000000010111111111111101111000000000000001100000000000011010000000000001111111111111111011111111111111001001111111111110111000000000000100000000000000010100000000000001110000000000000110000000000000001100000000000000010111111111101001000000000000000000000000000100000111111111100111011111111111010011111111111110111111111111110010111111111111000000000000000100001111111111101001111111111111100100000000000000010111111111111000111111111111110001111111111101000111111111110110100000000000011001111111111101010111111111111111000000000000111100000000000000001000000000010011011111111111010000000000000010100000000000000001011111111111110110000000000001100111111111111010011111111111101010000000000101100111111111110011011111111111000010000000000000011111111111111100100000000000011101111111111111100000000000000100100000000000100100000000000111000111111111110100111111111111111000000000000011100111111111101101000000000000010010000000000011001111111111110100100000000000000000000000000000000000000000000111100000000001000010000000000010001111111111111110100000000000011110000000000000100000000000000101000000000000000000000000000001010111111111110111100000000000000011111111111111111000000000001110100000000000101011111111111100000111111111111011011111111111110100000000000010111000000000001001100000000000001010000000000000001111111111111010100000000001100110000000000110001000000000001011100000000000000111111111111101011111111111101101111111111111111010000000000000111111111111110100111111111111010110000000000000011000000000000001111111111111111000000000000000011000000000001011000000000000111010000000000011011000000000010111000000000001100011111111111111110111111111111100000000000000011000000000000001010000000000000001111111111110111111111111111111111000000000000101100000000000011000000000000000100000000000001100111111111111100000000000000001001111111111111010111111111111111001111111111111010000000000000000100000000000001101111111111101011000000000000000000000000000010100000000000100011111111111110101011111111111111110000000000000111111111111101010011111111111001100000000000001111111111111111000011111111111111011111111111011001111111111110111011111111111100101111111111101101111111111111001100000000000010000000000000001100000000000000010111111111111111001111111111101001111111111110110000000000000011111111111111100110111111111110100100000000000000010000000000110101000000000001001011111111111011011111111111111110111111111111101100000000000101111111111111100101111111111111110100000000000011010000000000000100111111111111100100000000001011000000000000010100111111111111000000000000000000100000000000001101111111111111001100000000001000010000000000000111000000000000100100000000000010010000000000001010111111111100110111111111111111000000000000010110111111111101001100000000000010100000000000010011111111111111011011111111111010011111111111100111111111111110011011111111111111010000000000001101000000000001010111111111111011111111111111101001111111111110110000000000000001110000000000110001000000000000011111111111111010011111111111110101000000000000101000000000000101000000000000001010000000000000010000000000000001100000000000001010000000000000101100000000000011001111111111110010111111111111100111111111111100000000000000000000111111111111010011111111110110101111111111111110000000000000110011111111111101101111111111111011111111111100001111111111111001101111111111001010000000000000011100000000000000111111111111100011111111111110011000000000000011100000000000110100000000000001000100000000001001000000000000011001000000000000111100000000000000010000000000010011000000000001001000000000000000000000000000001101111111111111110111111111111011110000000000000101000000000000110100000000000001011111111111011010000000000000000000000000000010011111111111100110000000000001000100000000000001000000000000011011000000000000010011111111111100010000000000001101000000000000010111111111111111111111111111111011000000000000111011111111111111100000000000001010000000000001101011111111111100101111111111110101111111111111110011111111111010011111111111111010000000000000101000000000000001001111111111100110000000000000001100000000000000000000000000001101000000000000011100000000000001101111111111110110000000000001101100000000000100110000000000000000000000000001101000000000000101100000000000010101111111111110111011111111111010111111111111110011000000000000000011111111110100101111111111000010111111111111101011111111111000110000000000001111000000000000011100000000000110100000000000000110000000000001111000000000010001100000000000000010111111111111001011111111111110110000000000001101111111111111101100000000000011001111111111111010000000000000000011111111111110010000000000001100000000000001100011111111111111100000000000010101111111111111011100000000000010011111111111010111000000000100101100000000000101001111111111010110111111111111000111111111111101101111111111111011000000000000001111111111111110010000000000011111111111111111011011111111111100100000000000101000000000000000000000000000001001110000000000000110000000000000001100000000000111000000000000011000000000000000001100000000000010000000000000000110111111111111010100000000000010101111111111111011000000000000111111111111111001011111111111110001000000000000010111111111111101101111111111101010111111111110001111111111111011110000000000000101000000000000000100000000000001110000000000100000000000000000011111111111111101010000000000001001000000000000110100000000000001100000000000001111000000000001101011111111110110011111111111110101000000000011000011111111111101111111111111011010000000000001100011111111111010101111111111111101000000000001101000000000000000001111111111100010000000000001011000000000001001000000000000011000000000000001111000000000000001110000000000101100000000000010001100000000000100101111111111101111111111111111100111111111111010111111111111110000000000000000101100000000000010100000000000000011111111111111101000000000000101011111111111111100111111111111101000000000000000101111111111110110000000000000000000000000000000110000000000001000111111111111001011111111111111010000000000001000000000000000101011111111111011111111111111101111000000000001010000000000000111110000000000000001000000000000100111111111111111101111111111111101111111111111000011111111111011011111111111111010111111111111001111111111111101110000000000001101000000000000101111111111111110111111111111110110000000000000000011111111111001000000000000001100111111111110110011111111111011000000000000000010000000000000011100000000000101100000000000011011111111111111011111111111111100001111111111110101000000000000100011111111111111100000000000010001000000000000010000000000000010010000000000001001000000000000000000000000000001011111111111111100000000000000011011111111111011010000000000010001000000000001011000000000000010111111111111110000000000000000000011111111111000111111111111100111000000000001001111111111111001111111111111101111000000000000010000000000000000001111111111101000000000000010111100000000000001001111111111111001111111111110111011111111111001001111111111110110000000000000001011111111111101110000000000000001000000000001100000000000000010000000000000001101111111111111001111111111111100010000000000011010000000000001001111111111111111110000000000010001111111111111100111111111111101001111111111101111111111111111101100000000000101110000000000111001000000000000110011111111111011001111111111111111111111111110110011111111111100010000000000000010000000000000001000000000000101001111111111111110000000000001011111111111111100110000000000011101111111111111111011111111111010111111111111111001000000000010010011111111111011101111111111010100000000000000011111111111111010110000000000011011111111111111001111111111111011011111111111011010000000000000001000000000000000000000000000000001111111111111011011111111111100100000000000111010111111111110110011111111110101110000000000000100000000000001100011111111111111011111111111110010000000000000010111111111111110001111111110111110000000000000000000000000000001001111111111010100111111111110011011111111111011100000000000001011111111111111110011111111111101001111111111111100111111111111010011111111111001111111111111111001111111111101101100000000000001111111111111111110000000000010000000000000000001000000000000001011111111111110100011111111110100111111111110110100000000000000011100000000000010001111111111100101111111111111110100000000000011010000000000001101000000000000101100000000000000011111111111101110111111111110010011111111111101111111111111100000000000000010011000000000000100011111111111110011000000000001010011111111111000101111111111111110000000000001010100000000000010000000000000101010000000000000111011111111110110100000000000001101111111111110000011111111111100001111111111100010000000000010011111111111111111101111111111010100000000000001010111111111111100110000000000001011000000000000001000000000000111110000000000001110000000000100101000000000000011010000000000010010000000000001101111111111111010011111111111111001111111111110010011111111111100110000000000011000111111111111001000000000000111110000000000000100000000000001001011111111111110110000000000011101111111111110011100000000000000011111111110110000000000000001010111111111111101101111111111110110000000000000011100000000000010110000000000000000000000000000111000000000000000011111111111101001000000000000000011111111111101010000000000010110111111111111000000000000000010010000000000001011000000000000000111111111111101000000000000001100111111111111010011111111111110011111111111111111000000000000100000000000000011010000000000011100000000000000111000000000000010000000000000001000000000000001100111111111111100101111111111101001111111111111101100000000000010101111111111111001000000000000010100000000000010110000000000001100000000000000111111111111111110101111111111010111111111111111110011111111111001000000000000001111111111111101011111111111111100101111111111111100111111111111101000000000000000000000000000010110111111111111000011111111111001101111111111111000000000000001011011111111111010011111111111110100000000000000010100000000000110100000000000011010000000000001001111111111111100001111111111110000000000000000010100000000000010111111111111100011000000000001001011111111111101111111111111010001000000000000000000000000000011100000000000100011000000000001000000000000001000000000000000011001111111111110011111111111111110101111111111111001000000000000100100000000001000000000000000010110111111111111001111111111111110001111111111101110;
endcase
end
endmodule



module lut_weights_8(sbyte,addr);
input [3:0] addr;
output reg [20735:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b1000: sbyte = 20736'b000000000001001111111111111110101111111111101011000000000000110100000000000100111111111111011111111111111111011011111111101110000000000000000011000000000011000011111111111100100000000000010110111111111111101100000000000010000000000000001010000000000010001000000000000110011111111111001111000000000000111000000000001010101111111111100110111111111111001111111111110111000000000000010011111111111111101100000000000100111111111111001011000000000010101100000000000101100000000000100010111111111011100011111111110000101111111111100100111111111110111100000000000001110000000000001000000000000000000000000000000110000000000000000100000000000010110111111111101111001111111111101011000000000001011111111111111011000000000000000100111111111111000111111111111111001111111111110011000000000010100111111111111101110000000000000111111111111111101000000000000010111111111111100010111111111001011100000000000010111111111111111111111111111110010111111111111101111111111111110000111111111110111100000000000111101111111111110110000000000011001011111111110111011111111111011110111111111101111000000000001000110000000000011001111111111010111011111111111010100000000000101000000000000001101000000000000010010000000000010110000000000101010000000000000100110000000000000010111111111111111111111111111000010000000000101101111111111110011100000000000010011111111111001000000000000001101000000000000010110000000000000000000000000000011111111111111011011111111111011011111111111101101111111111111000100000000000001000111111111100111011111111111110000000000000010100111111111111001000000000000000001111111111111100111111111110001011111111111100110000000000011110111111111101101011111111101101010000000000100111111111111110110011111111110110000000000000010110000000000010000011111111111111100000000001000010000000000001111000000000001111001111111111011010111111111111000011111111110011010000000000101000000000000001011100000000000000010000000000100000000000000010011011111111110011100000000000001011111111111110000011111111110000000000000000100101111111111111110111111111110111011111111111110110111111111001110111111111110110011111111111110100111111111111101100000000001100100000000000000110111111111110001100000000000101011111111111111011111111111100100111111111101101001111111111101001111111111110001100000000000011100000000000010110111111111100110000000000000001110000000000000000000000000000011100000000001100100000000000100011111111111101110011111111111110000000000000010100000000000001011100000000000111101111111111100101000000000001001000000000001101001111111111010100111111111110000100000000000010000000000001000111000000000001010000000000000100000000000000010101111111111010111000000000010000111111111111111000111111111111101111111111110110100000000000000101111111111111011100000000000000110000000000110001111111111110110100000000001010111111111111110101000000000001001000000000000001000000000000000000111111111110110100000000000100011111111111100101000000000010001111111111111001110000000000101111000000000001111111111111111100111111111111111110111111111100110100000000000110110000000000100110000000000001100111111111111111001111111111111010000000000000011111111111111010110000000000001001000000000000101011111111111101001111111111011000111111111111110100000000000010110000000000001101111111111110101011111111111101101111111111100111111111111110010111111111111110010000000000011111111111111111010111111111110101111111111111111110111111111111111111111111110100100000000000000000111111111111101111111111111110100000000000001110111111111110100011111111111010010000000000101000000000000000110011111111111110000000000000010011111111111110111000000000010011110000000000100111111111111111101100000000010011011111111111101110000000000000101100000000010010110000000000001100111111111110100100000000001000010000000000000001000000000011011100000000000001011111111111111111000000000100011100000000010010100000000000111101111111111101111011111111111011101111111111010111111111111101101111111111101110011111111111100000111111111101101011111111111101011111111111011000111111111110001100000000001000110000000000101001000000000000001111111111110000101111111111101000000000000100001000000000000000001111111111011110111111111011110100000000000100010000000000010111000000000001111011111111111100000000000000000001111111111101010011111111110000100000000000001001000000000000000011111111111011110000000001001100111111111101111100000000000011110000000000001001111111111000100100000000000001100000000000001111111111111101111100000000001001000000000000100010000000000010011000000000000111011111111111011001000000000011100100000000000110100000000000011001111111111101010011111111111100100000000000000000000000000001010100000000001110110000000000000111000000000000101111111111101110111111111111110101111111111111011011111111111011010000000000000000111111111100000011111111111000100000000000011100000000000000010111111111111000000000000000000000111111111111010011111111111010011111111111101011111111111111001011111111111110101111111111100110111111111111110100000000011100000000000000110011111111111101111011111111110010111111111111011010000000000011100111111111110111111111111111000100000000000001100000000000001111010000000000011110111111111101010011111111111111011111111111010010000000000000110111111111111110011111111111111110111111111101111111111111110010001111111111010000000000000000011100000000001010100000000000010111111111111110011011111111111010011111111111010111000000000000000011111111111001000000000000001110111111111111110011111111111110100000000000000110111111111110010111111111111001101111111111001111000000000001111111111111110111110000000000011001111111111100111100000000000100001111111111101010000000000010111011111111111101111111111111101000111111111101111100000000001001111111111111111000111111111111010100000000000001101111111111011100111111111110011000000000000101000000000000011010000000000011101000000000000001001111111111001011000000000010000111111111111111011111111111110110000000000010000111111111110110111111111111111110111111111100010111111111111110100000000001001100000000000000010100000000000110100000000000111001111111111111010000000000001001100000000000100000111111111101110111111111111001010000000000001011111111111111111011111111101111010000000001010001000000000010000011111111110110101111111111110110111111111111111100000000001001111111111111111001000000000001011000000000001101000000000000111110111111111111011011111111111101111111111111111011000000000000011111111111111111011111111111111111111111111101110000000000001001011111111111110110111111111111100100000000000001110000000000011100111111111101110011111111110101101111111111101001000000000010010000000000000101001111111110101010111111111111101011111111111010101111111110111111111111111111011100000000010011010000000000011001000000000010101011111111111011011111111111100101000000000000101100000000000110110000000000011110000000000001011111111111111011100000000000000001111111111110101111111111110100101111111111011100111111111111101000000000000010001111111110111010000000000001000011111111101110010000000000000011111111111101100100000000010000100000000000011100111111111110011111111111111111010000000000010101111111111110011100000000000010100000000000001110111111111111101011111111111011110000000000110110000000000001111111111111111101110000000000001100000000000001010000000000000100110000000000001000000000000000010100000000000111001111111111110010000000000000010011111111111111011111111111011110111111111111000011111111110000110000000000000110111111111101010000000000001000100000000000010110111111111011101011111111111111110000000000001100111111111101000000000000000011100000000000000100000000000111000100000000000010000000000000101100000000000010011100000000000100001111111110111100000000000100001111111111100101111111111111000110000000000000110011111111111011011111111111110001111111111101001111111111111010101111111111100111111111111101111100000000000000101111111111110101000000000001110011111111111111111111111111110110111111111111011000000000010001010000000000000110111111111110011011111111111011010000000000111000000000000001100111111111110000111111111111110001000000000010111100000000010010111111111111010001000000000000011100000000000101000000000000001100000000000101110011111111111000101111111111110010111111111010000100000000001100001111111111011011000000000000101000000000000101110000000000110011000000000000000011111111110011011111111110110001000000000000011100000000010001000000000000000111111111111111110100000000001011011111111111111011111111111111010100000000001011011111111111110011000000000001000100000000001111101111111111100101000000000101100000000000001110001111111111010101111111111111110111111111111111101111111111111111111111111110111111111111111101101111111111010110111111111110000100000000010011000000000000010101111111111101011100000000000110011111111111101100000000000001011100000000000001011111111111001111000000000010101100000000010011101111111111010111000000000000010000000000010001100000000000001111111111111111101000000000001000000000000000000011000000000100000100000000001101111111111111110101111111111101101111111111111111000000000000000100111111111101011011111111111111101111111111011110000000000000000011111111110000000000000000000010000000000000111100000000000100010000000001000000111111111101001100000000000100111111111111000101000000000001000000000000010000110000000000000101000000000001010111111111111101110000000000000000111111111111101111111111111110001111111111111001111111111010011100000000000101110000000000000110111111111111001100000000000110011111111111101010111111111101110011111111111000100000000000011100111111111010111011111111111000011111111111000111000000000100110011111111110100010000000000100110111111111110111000000000000010100000000000001010111111111100100000000000000010000000000000011011000000000011011000000000000100000000000001011110111111111101111000000000010111001111111111100011111111111111100100000000000000001111111111110111111111111110111100000000001100011111111111110101000000000000000011111111110001001111111111101010111111111100111111111111111110011111111111100100000000000000101100000000000000101111111111101110111111111100011011111111111011000000000000010111000000000001000011111111111100010000000000000110000000000010010111111111111000001111111111110010000000000000100100000000001000111111111111110100000000000001101011111111111101001111111111111011000000000001100011111111111011010000000000111101000000000010111111111111111011000000000000100100000000000011010011111111111110100000000000001100111111111100001011111111111110000000000000101101000000000001010111111111111000010000000000100110000000000001000111111111110110101111111111000001000000000010011111111111111111011111111111101001000000000000000011111111111011011111111111110100111111111111111100000000000101010000000000110001000000000011000011111111101110011111111111100110000000000000010100000000000101000000000000100011111111111110010111111111111110100000000000111110111111111111110100000000000100110000000000010000111111111111110000000000000100010000000000000001000000000011111100000000001010001111111111100001111111111111101000000000000110111111111111111111000000000000111011111111111000010000000001001101111111111101001111111111110110011111111111101011111111111110011000000000010110011111111111110110111111111101100111111111110101100000000000001101111111111110011111111111110000011111111111111001000000000001101111111111101001000000000000111011000000000000000011111111110111010000000001100010111111111110100100000000001100000000000000111110000000000000100100000000000000001111111110110110000000000001011011111111101110000000000000100100111111111111010000000000001000100000000000010000111111111111110011111111111011100000000000000100000000000000110111111111110110100000000001000010000000000000000011111111111100001111111111010111000000000011101011111111111100101111111111001101111111111101011111111111111011100000000000010111111111111111011100000000000001011111111111001011111111111110101111111111111001110000000000011110000000000001111100000000001001010000000001000111111111111011010011111111111111110000000000001100111111111000010011111111111001111111111111101010111111111110101000000000000011010000000000100011000000000011110011111111110011101111111111110110111111111101100000000000001110110000000000001000000000000000011000000000000000100000000000010110111111111110001000000000000110001111111111000011000000000100011011111111111110010000000000110100000000000100010100000000000101101111111111000110000000000011000000000000001010000000000001001001000000000011001011111111111000100000000000100110000000000001011111111111110101010000000000010101111111111011101111111111111010010000000000010110111111111110111000000000000100110000000000101100000000000000111011111111111011101111111111100000111111111101011100000000000110111111111111001101000000000011100100000000000011110000000000011101000000000011000111111111100111101111111111110100111111111110111111111111111001010000000000001101111111111111010000000000001101100000000000101110000000000000000000000000000001010000000000101011000000000000111100000000000101011111111111011100111111111010111000000000001011001111111111001010111111111101110100000000001011111111111111011111000000000001100000000000001111111111111111100100000000000000010111111111111111100000000000011000000000000000000111111111111111010000000000000100111111111100111011111111110100111111111111100001111111111101011111111111111011110000000000110110111111111110001011111111111010001111111111111000000000000001111011111111110000000000000000111001111111111111011100000000000011111111111111111010111111111110000011111111110010001111111111101110000000000001000000000000000100100000000000110111111111111111000011111111111011110000000000010101111111111111110111111111111111100000000000100111111111111110110000000000000000001111111111101000000000000000100000000000001110100000000000000110000000000001001000000000000110000000000000000110000000000000010000000000001110010000000000101011000000000001100111111111110111110000000000100001000000000100101100000000001011000000000000110000000000000000001011111111111010111111111111001110000000000010101100000000000111011111111111101011111111111111100011111111111000101111111111100100111111111110101000000000000101110000000000011101111111111101111000000000000000001111111111100111111111111111110011111111111111001111111111101010111111111001101011111111101110110000000000001110000000000000000000000000001011111111111111010001111111111110111000000000000101100000000000110000000000000001010000000000000110100000000000111101000000000100011011111111111100110000000001000111111111111110011100000000000001101111111111101000111111111010110011111111111101101111111111101000000000000010000011111111111101101111111111100000000000000100010111111111111111000000000000000010111111111011111000000000001101100000000000101100111111111111110111111111110101000000000000011000111111111111101011111111111001100000000000011100111111111110011011111111110011100000000000111111111111111111110100000000001101101111111111111010000000000000100111111111101100101111111111011110000000000001011000000000001000110000000000110000111111111111001100000000010001001111111111000100000000000000101000000000000110101111111111001110000000000000011011111111110100101111111111000110111111111110110000000000010011110000000001100001000000000011100111111111111011101111111111111110111111111111111100000000000000001111111111101011000000000001111000000000000101111111111111110000111111111111110011111111101111110000000000100000111111111011011011111111111000001111111111011010111111111011110111111111110011110000000000011000111111111110110000000000000000110000000000100011111111111110010100000000000101000000000000110111000000000000111111111111111011010000000000000100111111111111111100000000001011111111111110011000111111111111001000000000001000111111111111111001000000000010101011111111101110110000000000110010000000000011110100000000001010011111111111010001111111111111011000000000000011111111111111111010000000000100010100000000001010100000000000010010111111111011101000000000000001011111111111100011111111111110111111111111110010100000000000111111111111111100100011111111111000001111111111010110111111111100101111111111110110001111111110011011111111111111101000000000010101010000000000010110111111111101101100000000000010101111111111011011000000000000001011111111111100110000000000100011111111111001110100000000000001100000000000000010000000000100111111111111111000010000000000001010111111111100101100000000000101011111111111110010000000000011110111111111111010110000000000011011000000000110100011111111110100001111111111011010111111111111010000000000001001110000000000000110000000000001111011111111110011101111111111001101000000000011111011111111111011011111111111111000000000000000001111111111111010000000000000000000111111111110011011111111111101001111111111110101111111111111011000000000000000001111111111100101111111111111101111111111111000011111111111101000000000000001011111111111101110111111111111110011111111111111101100000000000000010000000001000010000000000000001000000000010000110000000000010001111111111101001011111111110100111111111111011111111111111111110111111111111011010000000000010001000000000001000011111111111100000000000000011000111111111101000000000000000100101111111111101000000000000000010111111111110101010000000000011111000000000011011100000000001000011111111111001001000000000010010100000000000101101111111110111111000000000000101011111111111011000000000000100001000000000000110100000000001001111111111111010100000000000100001011111111110010011111111111000100111111111111111000000000000010100000000000000011111111111111111011111111111000100000000000110001111111111011101100000000000001101111111110111011000000000000000100000000010001001111111111010010111111111111101000000000000011000000000000010010000000000100101000000000000101011111111111111111111111111100101100000000000000111111111111111011111111111100001011111111110111001111111111111010000000000000011100000000001001110000000000000010111111111111001011111111110101101111111111111011111111111110111100000000000000010000000000101010000000000010110111111111111111011111111111110111111111111111111000000000000101010000000000000100111111111101100111111111111000011111111111111001111111111100000111111111111011110000000000011101000000000011110011111111110110111111111110100111000000000000110000000000010101001111111111010111111111111101100011111111111010101111111111011000111111111110101000000000001001101111111111010100111111111111011011111111111000011111111111100101000000000001001100000000001010011111111111110001111111111101001011111111110100100000000000101100111111111110011111111111111110100000000000011010111111111000011000000000000001111111111111000101111111111110011100000000000010100000000000110011000000000010000100000000000111011111111111111011111111111011001111111111111101000000000000000110000000000010100000000000011000010000000000101001000000000001110000000000000001010000000001000100111111111101000000000000001001110000000000010111111111111111101100000000001000010000000000110000111111111100011100000000000110100000000000011000111111111110011100000000000000010000000000011011000000000010010111111111111111110000000000100000000000000010110100000000000100111111111111101011111111111110111011111111110111100000000000111011000000000001011000000000000111100000000000101101111111111101000000000000000111101111111110111101000000000000100111111111111101000000000000110010000000000001011000000000000000101111111111100011000000000000001111111111111010011111111111010101111111111101111011111111101111100000000001000000000000000011111011111111110100111111111111110001111111111111010000000000000111010000000000000101000000000000100100000000000001011111111111011000000000000000100100000000000001011111111111101011111111111111110011111111111001110000000000010000111111111110111011111111111100001111111111111111111111111101100000000000000111011111111110110111111111111110001111111111111001101111111111011011111111111100011000000000001000010000000000001111000000000011011100000000010000011111111111100000000000000001011111111111111001001111111111000111111111111110110100000000001000011111111111101001111111111111111011111111111011110000000000010001000000000000110000000000000100000000000000100111111111111111001111111111101101011111111111001101000000000011011100000000001111010000000000011011111111111111000011111111111000101111111110110101111111111011011111111111111111010000000000101010111111111111000100000000001110010000000000001110111111111111111100000000000010011111111111111000000000000001010011111111110110100000000000011011000000000000100111111111111001010000000000000110111111111100111011111111111101011111111111110001111111111110000111111111111110011111111111100001;
endcase
end
endmodule



module lut_weights_9(sbyte,addr);
input [3:0] addr;
output reg [5759:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b1001: sbyte = 5760'b111111111100111111111111111100001111111111100000000000000011111011111111110100111111111111100110000000000010111011111111111111010000000010100010111111111101001011111111111100010000000000111100111111111110111011111111111001111111111111111011111111111001101100000000000100110000000000100100000000000101100011111111101110100000000000000111000000000100001011111111101000110000000000010110000000000001001000000000010000011111111111110111111111111000110011111111111111111111111111100101111111111000010011111111110100001111111111010010000000000000100100000000000101001111111111111100111111111111001000000000000000101111111111100110111111111111010100000000001010111111111111111011111111111101111111111111101101110000000000000011000000000100101111111111111011110000000000001111000000000001101011111111110010010000000000100010000000000000010100000000001001000000000000010001111111111010011011111111111001011111111110101000111111111110111111111111110011001111111111101000111111111101111011111111110110011111111111111101000000000001001100000000110000011111111111100101111111111011101000000000010010111111111111011000000000000011100100000000000000100000000000010110000000000000001100000000001001101111111111111001111111111101011100000000000101010000000000100011111111111101111111111111111100001111111111011001000000000011100111111111111101001111111111111101000000000001100100000000011011011111111111101011111111111101111000000000001001111111111111001001111111111101101011111111110011010000000000110110000000000001100111111111100100010000000000100110000000000101101000000000100010011111111111010011000000000111101111111111110011000000000000101110000000000001000011111111111110100000000001000101000000000100111000000000000111011111111111000101111111111101010000000000010010101111111110111100111111111101101011111111110010011111111111001000111111111110011100000000001000101111111111110011111111111101011000000000001100110000000000011100000000000000010011111111110101111111111111001000111111111110001100000000010000101111111111011111000000000100010000000000100110100000000001101001000000000011100111111111100101010000000000011011000000000011010100000000001010100000000000100000111111111100101100000000001111111111111111110111111111111101011011111111110000010000000001011001000000000000001111111111111010110000000000011100000000000000111000000000000100010000000000100110000000000011000111111111101110101111111111010111000000001000101111111111110101111111111111011011111111111100000111111111110100001111111110111000000000000010110111111111110110011111111111001110000000000001001111111111110010101111111111110110000000000001100111111111110100101111111110101111000000001001010011111111110100110000000000011000000000000001010100000000000010000000000001011011000000000011100100000000001100010000000000010100111111111101011000000000001010011111111111101011000000000001110100000000000000111111111111101111000000000011101100000000010001000000000001100111000000000110011111111111111000000000000000000100111111111100010000000000000001001111111111101100000000000010010111111111111000100000000000000101000000000010100100000000001010011111111110000010111111111111010011111111101110111111111111001001000000000101101000000000001101010000000001111000000000000001000100000000000101000000000000011110000000000111000000000000001100111111111111011010111111111110000000000000010111000000000000100111000000000000101100000000100000001111111110101110000000000001011111111111101010100000000000000011111111111111111100000000000011001111111111100010111111111100110111111111110000110000000000000100111111111011011000000000011011101111111111110010111111111110011111111111111111001111111111000111000000000010110111111111101000111111111110010110111111111010001011111111111100001111111111100101111111111111001011111111111110000000000000000000000000000000100100000000000100010000000000001111111111111100111111111111111000110000000010010111000000000010101011111111111011010000000000111001000000000010110111111111110110010000000001110011111111111100000011111111110101011111111111001100111111111111001000000000000000110000000000010101111111111111000000000000001010110000000000001100000000000010110111111111110010111111111111101010000000000100000000000000010011001111111111010101111111111111011000000000000010011111111110110001111111111111100011111111111000010000000000001110000000000000000000000000001011000000000000000000000000000011010100000000000011000000000001011001111111111101101011111111111110100000000000110010111111111110000011111111110111000000000000011001111111111101100011111111110110101111111111101000000000000100111111111111111010000000000001011001000000000011010111111111101101101111111111111010000000000010001011111111111101100000000001001000111111111110000100000000010011101111111111011111111111111110000111111111101100000000000001010101000000000001011000000000010000001111111110011000111111111101001100000000010110010000000001100111000000000101001000000000010111111111111111011110111111111101100000000000000111101111111111010011000000000010000011111111110101111111111111100110000000000010011011111111111101111111111111100101000000000001100111111111111001101111111111100010000000000100000100000000000011011111111111110001000000000010100011111111111100110000000000000000000000000000111111111111111011101111111111101110000000001000101011111111111000001111111111111011111111111101000011111111101111101111111111111000111111111011011111111111110101001111111111010010000000000111100011111111110111000000000000010110000000000000001111111111111011011111111111010101111111111101100100000000000111011111111111010111000000000100111100000000000100010000000001110010111111111100110111111111111000010000000000010010111111111101000100000000000100011111111111010111000000000010001111111111111010101111111111011010;
endcase
end
endmodule



