module lut_biases_1(sbyte,addr);
input [3:0] addr;
output reg [191:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0001: sbyte = 192'b000000000000000100000000011111010000000000100111000000000000001111111111111100000000000000000001000000000100000111111111111001000000000001100100000000000011000100000000000110110000000001000100;
endcase
end
endmodule



module lut_biases_2(sbyte,addr);
input [3:0] addr;
output reg [191:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0010: sbyte = 192'b000000000000010100000000000111010000000000110000000000000000000011111111111101010000000000011100000000000000000000000000000011110000000000100111000000000001001000000000000001001111111111110010;
endcase
end
endmodule



module lut_biases_3(sbyte,addr);
input [3:0] addr;
output reg [191:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0011: sbyte = 192'b000000000001101011111111111100100000000000000000000000000001100011111111111101010000000000000000000000000000100100000000000101010000000000101110000000000010110000000000000011111111111111110100;
endcase
end
endmodule



module lut_biases_4(sbyte,addr);
input [3:0] addr;
output reg [383:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0100: sbyte = 384'b111111111111101000000000000000110000000000111111000000000000110011111111111101000000000000010111000000000001110011111111111101101111111111111001000000000011010111111111111110000000000000000011000000000010110000000000000011010000000000001111111111111111101100000000000000110000000000011101111111111111101100000000000100000000000000001010000000000001001011111111111011011111111111111000;
endcase
end
endmodule



module lut_biases_5(sbyte,addr);
input [3:0] addr;
output reg [383:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0101: sbyte = 384'b000000000000111100000000000001001111111111111100000000000001000100000000000101100000000000001101000000000000100011111111111110110000000000000101111111111111110011111111111111100000000000000000000000000010011100000000000110101111111111111101111111111111111100000000000001110000000000000000000000000001100100000000000011101111111111110110111111111111010011111111111111000000000000010010;
endcase
end
endmodule



module lut_biases_6(sbyte,addr);
input [3:0] addr;
output reg [383:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0110: sbyte = 384'b111111111111100000000000000101000000000000001111000000000000000000000000000000011111111111110100000000000000111011111111111111100000000000001110000000000000001100000000000101010000000000000000000000000000001011111111111111110000000000001010000000000001001000000000000000111111111111111011111111111111110100000000000001010000000000000000000000000000100000000000000001100000000000000111;
endcase
end
endmodule



module lut_biases_7(sbyte,addr);
input [3:0] addr;
output reg [575:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0111: sbyte = 576'b000000000000001111111111111110000000000000010111000000000000100000000000000000011111111111101011111111111111010100000000000001011111111111111011111111111111111111111111111100010000000000000011000000000001001111111111111100111111111111111101111111111111110111111111111100111111111111111000000000000000000011111111111111100000000000000101000000000000100100000000000000010000000000000101000000000000010100000000000011101111111111110010000000000000000000000000000010101111111111111101111111111111111100000000000101001111111111110101000000000000000000000000000100010000000000000110;
endcase
end
endmodule



module lut_biases_8(sbyte,addr);
input [3:0] addr;
output reg [575:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b1000: sbyte = 576'b000000000000111111111111111011100000000000000001111111111111010111111111111111101111111111100110111111111111101000000000000110101111111111111101111111111110100111111111111010100000000000000111111111111111000100000000000100100000000000000010000000000001011100000000000000001111111111111110000000000001000000000000000000100000000000011111000000000000100100000000001111111111111111101101111111111111110111111111111011111111111111101001111111111111111111111111111111101111111111110011111111111111110000000000000000111111111111110001000000000000100111111111111111100000000000010100;
endcase
end
endmodule



module lut_biases_9(sbyte,addr);
input [3:0] addr;
output reg [159:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b1001: sbyte = 160'b1111111111110000111111111111011111111111110111011111111111100000111111111110101000000000001100100000000000000101000000000000011000000000000101101111111111110010;
endcase
end
endmodule



