module lut_index_1(sbyte,addr);
input [3:0] addr;
output reg [26:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0001: sbyte = 27'b000000000000000000000000000;
endcase
end
endmodule



module lut_index_2(sbyte,addr);
input [3:0] addr;
output reg [323:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0010: sbyte = 324'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endcase
end
endmodule



module lut_index_3(sbyte,addr);
input [3:0] addr;
output reg [323:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0011: sbyte = 324'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endcase
end
endmodule



module lut_index_4(sbyte,addr);
input [3:0] addr;
output reg [323:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0100: sbyte = 324'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endcase
end
endmodule



module lut_index_5(sbyte,addr);
input [3:0] addr;
output reg [647:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0101: sbyte = 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endcase
end
endmodule



module lut_index_6(sbyte,addr);
input [3:0] addr;
output reg [647:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0110: sbyte = 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endcase
end
endmodule



module lut_index_7(sbyte,addr);
input [3:0] addr;
output reg [647:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b0111: sbyte = 648'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endcase
end
endmodule



module lut_index_8(sbyte,addr);
input [3:0] addr;
output reg [107:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b1000: sbyte = 108'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endcase
end
endmodule



module lut_index_9(sbyte,addr);
input [3:0] addr;
output reg [107:0] sbyte;

always @ (addr) begin

(* synthesis, full_case, parallel_case *) case (addr)

4'b1001: sbyte = 108'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endcase
end
endmodule



